// This is the unpowered netlist.
module DSP (Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    Tile_X0Y0_E1BEG,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2BEG,
    Tile_X0Y0_E2BEGb,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6BEG,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4BEG,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_NN4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_SS4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W1END,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W2END,
    Tile_X0Y0_W2MID,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_W6END,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y0_WW4END,
    Tile_X0Y1_E1BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2BEG,
    Tile_X0Y1_E2BEGb,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6BEG,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4BEG,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_NN4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_SS4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W1END,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W2END,
    Tile_X0Y1_W2MID,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_W6END,
    Tile_X0Y1_WW4BEG,
    Tile_X0Y1_WW4END);
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output [3:0] Tile_X0Y0_E1BEG;
 input [3:0] Tile_X0Y0_E1END;
 output [7:0] Tile_X0Y0_E2BEG;
 output [7:0] Tile_X0Y0_E2BEGb;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 output [11:0] Tile_X0Y0_E6BEG;
 input [11:0] Tile_X0Y0_E6END;
 output [15:0] Tile_X0Y0_EE4BEG;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 output [15:0] Tile_X0Y0_NN4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 input [15:0] Tile_X0Y0_SS4END;
 output [3:0] Tile_X0Y0_W1BEG;
 input [3:0] Tile_X0Y0_W1END;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 input [7:0] Tile_X0Y0_W2END;
 input [7:0] Tile_X0Y0_W2MID;
 output [11:0] Tile_X0Y0_W6BEG;
 input [11:0] Tile_X0Y0_W6END;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [15:0] Tile_X0Y0_WW4END;
 output [3:0] Tile_X0Y1_E1BEG;
 input [3:0] Tile_X0Y1_E1END;
 output [7:0] Tile_X0Y1_E2BEG;
 output [7:0] Tile_X0Y1_E2BEGb;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 output [11:0] Tile_X0Y1_E6BEG;
 input [11:0] Tile_X0Y1_E6END;
 output [15:0] Tile_X0Y1_EE4BEG;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 input [15:0] Tile_X0Y1_NN4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [15:0] Tile_X0Y1_SS4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 input [3:0] Tile_X0Y1_W1END;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 input [7:0] Tile_X0Y1_W2END;
 input [7:0] Tile_X0Y1_W2MID;
 output [11:0] Tile_X0Y1_W6BEG;
 input [11:0] Tile_X0Y1_W6END;
 output [15:0] Tile_X0Y1_WW4BEG;
 input [15:0] Tile_X0Y1_WW4END;

 wire \Tile_X0Y0_DSP_top/ConfigBits[0] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[100] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[101] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[102] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[103] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[104] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[105] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[106] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[107] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[108] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[109] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[10] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[110] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[111] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[112] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[113] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[114] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[115] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[116] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[117] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[118] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[119] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[11] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[120] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[121] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[122] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[123] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[124] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[125] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[126] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[127] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[128] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[129] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[12] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[130] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[131] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[132] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[133] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[134] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[135] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[136] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[137] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[138] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[139] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[13] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[140] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[141] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[142] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[143] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[144] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[145] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[146] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[147] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[148] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[149] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[14] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[150] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[151] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[152] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[153] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[154] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[155] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[156] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[157] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[158] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[159] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[15] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[160] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[161] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[162] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[163] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[164] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[165] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[166] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[167] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[168] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[169] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[16] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[170] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[171] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[172] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[173] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[174] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[175] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[176] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[177] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[178] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[179] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[17] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[180] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[181] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[182] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[183] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[184] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[185] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[186] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[187] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[188] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[189] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[18] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[190] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[191] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[192] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[193] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[194] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[195] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[196] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[197] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[198] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[199] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[19] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[1] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[200] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[201] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[202] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[203] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[204] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[205] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[206] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[207] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[208] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[209] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[20] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[210] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[211] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[212] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[213] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[214] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[215] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[216] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[217] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[218] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[219] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[21] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[220] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[221] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[222] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[223] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[224] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[225] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[226] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[227] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[228] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[229] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[22] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[230] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[231] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[232] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[233] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[234] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[235] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[236] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[237] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[238] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[239] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[23] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[240] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[241] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[242] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[243] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[244] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[245] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[246] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[247] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[248] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[249] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[24] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[250] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[251] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[252] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[253] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[254] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[255] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[256] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[257] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[258] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[259] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[25] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[260] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[261] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[262] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[263] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[264] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[265] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[266] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[267] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[268] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[269] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[26] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[270] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[271] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[272] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[273] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[274] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[275] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[276] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[277] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[278] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[279] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[27] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[280] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[281] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[282] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[283] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[284] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[285] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[286] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[287] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[288] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[289] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[28] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[290] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[291] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[292] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[293] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[294] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[295] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[296] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[297] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[298] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[299] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[29] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[2] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[300] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[301] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[302] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[303] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[304] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[305] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[306] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[307] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[308] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[309] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[30] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[310] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[311] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[312] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[313] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[314] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[315] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[316] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[317] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[318] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[319] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[31] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[320] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[321] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[322] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[323] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[324] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[325] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[326] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[327] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[328] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[329] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[32] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[330] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[331] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[332] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[333] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[334] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[335] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[336] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[337] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[338] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[339] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[33] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[340] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[341] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[342] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[343] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[344] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[345] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[346] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[347] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[348] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[349] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[34] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[350] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[351] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[352] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[353] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[354] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[355] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[356] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[357] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[358] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[359] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[35] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[360] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[361] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[362] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[363] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[364] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[365] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[366] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[367] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[368] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[369] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[36] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[370] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[371] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[372] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[373] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[374] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[375] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[376] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[377] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[378] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[379] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[37] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[380] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[381] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[382] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[383] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[384] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[385] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[386] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[387] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[388] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[389] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[38] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[390] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[391] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[392] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[393] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[394] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[395] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[396] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[397] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[398] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[399] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[39] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[3] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[400] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[401] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[402] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[403] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[404] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[405] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[40] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[41] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[42] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[43] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[44] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[45] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[46] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[47] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[48] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[49] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[4] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[50] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[51] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[52] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[53] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[54] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[55] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[56] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[57] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[58] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[59] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[5] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[60] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[61] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[62] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[63] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[64] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[65] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[66] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[67] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[68] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[69] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[6] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[70] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[71] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[72] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[73] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[74] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[75] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[76] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[77] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[78] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[79] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[7] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[80] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[81] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[82] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[83] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[84] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[85] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[86] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[87] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[88] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[89] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[8] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[90] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[91] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[92] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[93] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[94] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[95] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[96] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[97] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[98] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[99] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits[9] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[0] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[100] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[101] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[102] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[103] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[104] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[105] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[106] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[107] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[108] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[109] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[10] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[110] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[111] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[112] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[113] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[114] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[115] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[116] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[117] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[118] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[119] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[11] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[120] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[121] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[122] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[123] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[124] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[125] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[126] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[127] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[128] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[129] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[12] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[130] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[131] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[132] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[133] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[134] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[135] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[136] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[137] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[138] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[139] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[13] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[140] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[141] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[142] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[143] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[144] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[145] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[146] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[147] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[148] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[149] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[14] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[150] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[151] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[152] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[153] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[154] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[155] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[156] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[157] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[158] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[159] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[15] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[160] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[161] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[162] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[163] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[164] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[165] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[166] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[167] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[168] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[169] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[16] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[170] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[171] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[172] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[173] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[174] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[175] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[176] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[177] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[178] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[179] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[17] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[180] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[181] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[182] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[183] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[184] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[185] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[186] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[187] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[188] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[189] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[18] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[190] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[191] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[192] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[193] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[194] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[195] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[196] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[197] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[198] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[199] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[19] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[1] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[200] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[201] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[202] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[203] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[204] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[205] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[206] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[207] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[208] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[209] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[20] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[210] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[211] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[212] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[213] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[214] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[215] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[216] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[217] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[218] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[219] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[21] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[220] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[221] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[222] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[223] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[224] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[225] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[226] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[227] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[228] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[229] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[22] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[230] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[231] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[232] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[233] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[234] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[235] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[236] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[237] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[238] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[239] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[23] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[240] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[241] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[242] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[243] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[244] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[245] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[246] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[247] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[248] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[249] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[24] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[250] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[251] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[252] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[253] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[254] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[255] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[256] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[257] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[258] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[259] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[25] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[260] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[261] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[262] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[263] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[264] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[265] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[266] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[267] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[268] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[269] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[26] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[270] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[271] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[272] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[273] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[274] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[275] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[276] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[277] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[278] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[279] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[27] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[280] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[281] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[282] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[283] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[284] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[285] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[286] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[287] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[288] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[289] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[28] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[290] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[291] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[292] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[293] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[294] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[295] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[296] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[297] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[298] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[299] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[29] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[2] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[300] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[301] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[302] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[303] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[304] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[305] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[306] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[307] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[308] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[309] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[30] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[310] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[311] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[312] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[313] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[314] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[315] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[316] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[317] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[318] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[319] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[31] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[320] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[321] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[322] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[323] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[324] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[325] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[326] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[327] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[328] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[329] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[32] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[330] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[331] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[332] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[333] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[334] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[335] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[336] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[337] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[338] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[339] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[33] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[340] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[341] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[342] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[343] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[344] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[345] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[346] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[347] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[348] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[349] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[34] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[350] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[351] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[352] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[353] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[354] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[355] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[356] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[357] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[358] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[359] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[35] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[360] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[361] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[362] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[363] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[364] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[365] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[366] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[367] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[368] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[369] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[36] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[370] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[371] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[372] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[373] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[374] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[375] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[376] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[377] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[378] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[379] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[37] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[380] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[381] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[382] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[383] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[384] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[385] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[386] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[387] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[388] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[389] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[38] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[390] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[391] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[392] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[393] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[394] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[395] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[396] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[397] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[398] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[399] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[39] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[3] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[400] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[401] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[402] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[403] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[404] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[405] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[40] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[41] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[42] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[43] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[44] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[45] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[46] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[47] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[48] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[49] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[4] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[50] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[51] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[52] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[53] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[54] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[55] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[56] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[57] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[58] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[59] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[5] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[60] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[61] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[62] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[63] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[64] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[65] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[66] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[67] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[68] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[69] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[6] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[70] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[71] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[72] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[73] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[74] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[75] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[76] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[77] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[78] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[79] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[7] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[80] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[81] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[82] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[83] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[84] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[85] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[86] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[87] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[88] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[89] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[8] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[90] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[91] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[92] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[93] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[94] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[95] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[96] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[97] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[98] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[99] ;
 wire \Tile_X0Y0_DSP_top/ConfigBits_N[9] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/E6BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/EE4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[0] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[10] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[11] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[12] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[13] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[14] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[15] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[16] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[17] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[18] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[19] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[1] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[20] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[21] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[22] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[23] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[24] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[25] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[26] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[27] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[28] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[29] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[2] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[30] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[31] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[3] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[4] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[5] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[6] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[7] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[8] ;
 wire \Tile_X0Y0_DSP_top/FrameData_O_i[9] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[0] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[10] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[11] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[12] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[13] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[14] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[15] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[16] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[17] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[18] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[19] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[1] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[2] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[3] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[4] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[5] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[6] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[7] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[8] ;
 wire \Tile_X0Y0_DSP_top/FrameStrobe_O_i[9] ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out0 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out1 ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_0_ ;
 wire \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_1_ ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_ABb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_EFb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHa_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J2MID_GHb_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JE2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JN2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JS2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[0] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[1] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[2] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[3] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[4] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[5] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[6] ;
 wire \Tile_X0Y0_DSP_top/JW2BEG[7] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_AB_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_CD_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_EF_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[0] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[1] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[2] ;
 wire \Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/N4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/NN4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/S4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/SS4BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/W6BEG_i[9] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[0] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[10] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[11] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[1] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[2] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[3] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[4] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[5] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[6] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[7] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[8] ;
 wire \Tile_X0Y0_DSP_top/WW4BEG_i[9] ;
 wire \Tile_X0Y0_S1BEG[0] ;
 wire \Tile_X0Y0_S1BEG[1] ;
 wire \Tile_X0Y0_S1BEG[2] ;
 wire \Tile_X0Y0_S1BEG[3] ;
 wire \Tile_X0Y0_S2BEG[0] ;
 wire \Tile_X0Y0_S2BEG[1] ;
 wire \Tile_X0Y0_S2BEG[2] ;
 wire \Tile_X0Y0_S2BEG[3] ;
 wire \Tile_X0Y0_S2BEG[4] ;
 wire \Tile_X0Y0_S2BEG[5] ;
 wire \Tile_X0Y0_S2BEG[6] ;
 wire \Tile_X0Y0_S2BEG[7] ;
 wire \Tile_X0Y0_S2BEGb[0] ;
 wire \Tile_X0Y0_S2BEGb[1] ;
 wire \Tile_X0Y0_S2BEGb[2] ;
 wire \Tile_X0Y0_S2BEGb[3] ;
 wire \Tile_X0Y0_S2BEGb[4] ;
 wire \Tile_X0Y0_S2BEGb[5] ;
 wire \Tile_X0Y0_S2BEGb[6] ;
 wire \Tile_X0Y0_S2BEGb[7] ;
 wire \Tile_X0Y0_S4BEG[0] ;
 wire \Tile_X0Y0_S4BEG[10] ;
 wire \Tile_X0Y0_S4BEG[11] ;
 wire \Tile_X0Y0_S4BEG[12] ;
 wire \Tile_X0Y0_S4BEG[13] ;
 wire \Tile_X0Y0_S4BEG[14] ;
 wire \Tile_X0Y0_S4BEG[15] ;
 wire \Tile_X0Y0_S4BEG[1] ;
 wire \Tile_X0Y0_S4BEG[2] ;
 wire \Tile_X0Y0_S4BEG[3] ;
 wire \Tile_X0Y0_S4BEG[4] ;
 wire \Tile_X0Y0_S4BEG[5] ;
 wire \Tile_X0Y0_S4BEG[6] ;
 wire \Tile_X0Y0_S4BEG[7] ;
 wire \Tile_X0Y0_S4BEG[8] ;
 wire \Tile_X0Y0_S4BEG[9] ;
 wire \Tile_X0Y0_SS4BEG[0] ;
 wire \Tile_X0Y0_SS4BEG[10] ;
 wire \Tile_X0Y0_SS4BEG[11] ;
 wire \Tile_X0Y0_SS4BEG[12] ;
 wire \Tile_X0Y0_SS4BEG[13] ;
 wire \Tile_X0Y0_SS4BEG[14] ;
 wire \Tile_X0Y0_SS4BEG[15] ;
 wire \Tile_X0Y0_SS4BEG[1] ;
 wire \Tile_X0Y0_SS4BEG[2] ;
 wire \Tile_X0Y0_SS4BEG[3] ;
 wire \Tile_X0Y0_SS4BEG[4] ;
 wire \Tile_X0Y0_SS4BEG[5] ;
 wire \Tile_X0Y0_SS4BEG[6] ;
 wire \Tile_X0Y0_SS4BEG[7] ;
 wire \Tile_X0Y0_SS4BEG[8] ;
 wire \Tile_X0Y0_SS4BEG[9] ;
 wire \Tile_X0Y0_top2bot[0] ;
 wire \Tile_X0Y0_top2bot[10] ;
 wire \Tile_X0Y0_top2bot[11] ;
 wire \Tile_X0Y0_top2bot[12] ;
 wire \Tile_X0Y0_top2bot[13] ;
 wire \Tile_X0Y0_top2bot[14] ;
 wire \Tile_X0Y0_top2bot[15] ;
 wire \Tile_X0Y0_top2bot[16] ;
 wire \Tile_X0Y0_top2bot[17] ;
 wire \Tile_X0Y0_top2bot[1] ;
 wire \Tile_X0Y0_top2bot[2] ;
 wire \Tile_X0Y0_top2bot[3] ;
 wire \Tile_X0Y0_top2bot[4] ;
 wire \Tile_X0Y0_top2bot[5] ;
 wire \Tile_X0Y0_top2bot[6] ;
 wire \Tile_X0Y0_top2bot[7] ;
 wire \Tile_X0Y0_top2bot[8] ;
 wire \Tile_X0Y0_top2bot[9] ;
 wire \Tile_X0Y1_DSP_bot/A0 ;
 wire \Tile_X0Y1_DSP_bot/A1 ;
 wire \Tile_X0Y1_DSP_bot/A2 ;
 wire \Tile_X0Y1_DSP_bot/A3 ;
 wire \Tile_X0Y1_DSP_bot/A4 ;
 wire \Tile_X0Y1_DSP_bot/A5 ;
 wire \Tile_X0Y1_DSP_bot/A6 ;
 wire \Tile_X0Y1_DSP_bot/A7 ;
 wire \Tile_X0Y1_DSP_bot/B0 ;
 wire \Tile_X0Y1_DSP_bot/B1 ;
 wire \Tile_X0Y1_DSP_bot/B2 ;
 wire \Tile_X0Y1_DSP_bot/B3 ;
 wire \Tile_X0Y1_DSP_bot/B4 ;
 wire \Tile_X0Y1_DSP_bot/B5 ;
 wire \Tile_X0Y1_DSP_bot/B6 ;
 wire \Tile_X0Y1_DSP_bot/B7 ;
 wire \Tile_X0Y1_DSP_bot/C0 ;
 wire \Tile_X0Y1_DSP_bot/C1 ;
 wire \Tile_X0Y1_DSP_bot/C10 ;
 wire \Tile_X0Y1_DSP_bot/C11 ;
 wire \Tile_X0Y1_DSP_bot/C12 ;
 wire \Tile_X0Y1_DSP_bot/C13 ;
 wire \Tile_X0Y1_DSP_bot/C14 ;
 wire \Tile_X0Y1_DSP_bot/C15 ;
 wire \Tile_X0Y1_DSP_bot/C16 ;
 wire \Tile_X0Y1_DSP_bot/C17 ;
 wire \Tile_X0Y1_DSP_bot/C18 ;
 wire \Tile_X0Y1_DSP_bot/C19 ;
 wire \Tile_X0Y1_DSP_bot/C2 ;
 wire \Tile_X0Y1_DSP_bot/C3 ;
 wire \Tile_X0Y1_DSP_bot/C4 ;
 wire \Tile_X0Y1_DSP_bot/C5 ;
 wire \Tile_X0Y1_DSP_bot/C6 ;
 wire \Tile_X0Y1_DSP_bot/C7 ;
 wire \Tile_X0Y1_DSP_bot/C8 ;
 wire \Tile_X0Y1_DSP_bot/C9 ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[0] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[100] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[101] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[102] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[103] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[104] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[105] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[106] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[107] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[108] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[109] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[10] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[110] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[111] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[112] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[113] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[114] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[115] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[116] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[117] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[118] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[119] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[11] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[120] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[121] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[122] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[123] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[124] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[125] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[126] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[127] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[128] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[129] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[12] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[130] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[131] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[132] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[133] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[134] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[135] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[136] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[137] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[138] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[139] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[13] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[140] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[141] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[142] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[143] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[144] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[145] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[146] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[147] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[148] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[149] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[14] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[150] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[151] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[152] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[153] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[154] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[155] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[156] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[157] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[158] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[159] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[15] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[160] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[161] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[162] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[163] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[164] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[165] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[166] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[167] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[168] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[169] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[16] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[170] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[171] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[172] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[173] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[174] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[175] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[176] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[177] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[178] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[179] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[17] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[180] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[181] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[182] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[183] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[184] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[185] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[186] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[187] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[188] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[189] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[18] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[190] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[191] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[192] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[193] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[194] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[195] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[196] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[197] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[198] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[199] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[19] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[1] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[200] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[201] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[202] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[203] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[204] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[205] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[206] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[207] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[208] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[209] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[20] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[210] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[211] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[212] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[213] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[214] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[215] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[216] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[217] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[218] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[219] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[21] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[220] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[221] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[222] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[223] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[224] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[225] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[226] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[227] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[228] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[229] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[22] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[230] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[231] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[232] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[233] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[234] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[235] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[236] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[237] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[238] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[239] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[23] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[240] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[241] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[242] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[243] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[244] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[245] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[246] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[247] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[248] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[249] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[24] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[250] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[251] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[252] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[253] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[254] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[255] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[256] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[257] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[258] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[259] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[25] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[260] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[261] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[262] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[263] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[264] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[265] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[266] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[267] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[268] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[269] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[26] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[270] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[271] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[272] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[273] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[274] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[275] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[276] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[277] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[278] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[279] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[27] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[280] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[281] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[282] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[283] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[284] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[285] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[286] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[287] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[288] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[289] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[28] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[290] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[291] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[292] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[293] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[294] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[295] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[296] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[297] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[298] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[299] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[29] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[2] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[300] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[301] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[302] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[303] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[304] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[305] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[306] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[307] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[308] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[309] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[30] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[310] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[311] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[312] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[313] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[314] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[315] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[316] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[317] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[318] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[319] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[31] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[320] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[321] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[322] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[323] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[324] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[325] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[326] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[327] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[328] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[329] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[32] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[330] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[331] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[332] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[333] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[334] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[335] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[336] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[337] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[338] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[339] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[33] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[340] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[341] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[342] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[343] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[344] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[345] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[346] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[347] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[348] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[349] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[34] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[350] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[351] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[352] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[353] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[354] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[355] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[356] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[357] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[358] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[359] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[35] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[360] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[361] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[362] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[363] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[364] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[365] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[366] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[367] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[368] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[369] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[36] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[370] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[371] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[372] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[373] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[374] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[375] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[376] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[377] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[378] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[379] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[37] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[380] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[381] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[382] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[383] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[384] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[385] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[386] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[387] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[388] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[389] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[38] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[390] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[391] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[392] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[393] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[394] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[395] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[396] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[397] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[398] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[399] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[39] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[3] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[400] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[401] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[402] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[403] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[404] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[405] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[406] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[407] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[408] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[409] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[40] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[410] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[411] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[412] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[413] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[414] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[415] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[41] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[42] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[43] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[44] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[45] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[46] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[47] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[48] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[49] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[4] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[50] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[51] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[52] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[53] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[54] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[55] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[56] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[57] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[58] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[59] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[5] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[60] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[61] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[62] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[63] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[64] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[65] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[66] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[67] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[68] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[69] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[6] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[70] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[71] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[72] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[73] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[74] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[75] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[76] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[77] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[78] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[79] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[7] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[80] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[81] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[82] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[83] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[84] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[85] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[86] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[87] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[88] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[89] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[8] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[90] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[91] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[92] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[93] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[94] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[95] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[96] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[97] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[98] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[99] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits[9] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[0] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[100] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[101] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[102] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[103] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[104] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[105] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[106] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[107] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[108] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[109] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[10] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[110] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[111] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[112] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[113] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[114] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[115] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[116] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[117] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[118] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[119] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[11] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[120] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[121] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[122] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[123] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[124] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[125] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[126] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[127] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[128] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[129] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[12] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[130] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[131] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[132] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[133] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[134] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[135] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[136] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[137] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[138] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[139] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[13] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[140] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[141] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[142] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[143] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[144] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[145] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[146] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[147] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[148] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[149] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[14] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[150] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[151] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[152] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[153] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[154] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[155] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[156] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[157] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[158] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[159] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[15] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[160] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[161] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[162] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[163] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[164] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[165] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[166] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[167] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[168] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[169] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[16] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[170] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[171] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[172] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[173] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[174] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[175] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[176] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[177] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[178] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[179] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[17] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[180] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[181] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[182] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[183] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[184] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[185] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[186] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[187] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[188] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[189] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[18] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[190] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[191] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[192] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[193] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[194] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[195] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[196] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[197] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[198] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[199] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[19] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[1] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[200] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[201] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[202] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[203] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[204] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[205] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[206] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[207] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[208] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[209] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[20] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[210] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[211] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[212] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[213] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[214] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[215] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[216] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[217] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[218] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[219] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[21] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[220] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[221] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[222] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[223] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[224] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[225] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[226] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[227] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[228] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[229] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[22] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[230] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[231] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[232] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[233] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[234] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[235] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[236] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[237] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[238] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[239] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[23] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[240] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[241] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[242] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[243] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[244] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[245] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[246] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[247] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[248] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[249] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[24] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[250] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[251] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[252] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[253] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[254] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[255] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[256] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[257] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[258] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[259] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[25] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[260] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[261] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[262] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[263] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[264] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[265] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[266] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[267] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[268] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[269] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[26] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[270] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[271] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[272] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[273] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[274] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[275] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[276] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[277] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[278] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[279] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[27] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[280] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[281] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[282] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[283] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[284] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[285] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[286] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[287] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[288] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[289] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[28] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[290] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[291] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[292] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[293] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[294] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[295] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[296] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[297] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[298] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[299] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[29] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[2] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[300] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[301] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[302] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[303] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[304] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[305] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[306] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[307] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[308] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[309] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[30] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[310] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[311] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[312] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[313] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[314] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[315] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[316] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[317] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[318] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[319] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[31] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[320] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[321] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[322] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[323] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[324] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[325] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[326] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[327] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[328] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[329] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[32] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[330] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[331] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[332] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[333] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[334] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[335] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[336] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[337] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[338] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[339] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[33] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[340] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[341] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[342] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[343] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[344] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[345] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[346] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[347] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[348] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[349] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[34] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[350] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[351] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[352] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[353] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[354] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[355] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[356] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[357] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[358] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[359] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[35] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[360] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[361] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[362] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[363] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[364] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[365] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[366] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[367] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[368] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[369] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[36] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[370] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[371] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[372] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[373] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[374] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[375] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[376] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[377] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[378] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[379] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[37] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[380] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[381] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[382] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[383] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[384] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[385] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[386] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[387] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[388] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[389] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[38] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[390] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[391] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[392] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[393] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[394] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[395] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[396] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[397] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[398] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[399] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[39] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[3] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[400] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[401] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[402] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[403] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[404] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[405] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[406] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[407] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[408] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[409] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[40] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[410] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[411] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[412] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[413] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[414] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[415] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[41] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[42] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[43] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[44] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[45] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[46] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[47] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[48] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[49] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[4] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[50] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[51] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[52] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[53] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[54] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[55] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[56] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[57] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[58] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[59] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[5] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[60] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[61] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[62] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[63] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[64] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[65] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[66] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[67] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[68] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[69] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[6] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[70] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[71] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[72] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[73] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[74] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[75] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[76] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[77] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[78] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[79] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[7] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[80] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[81] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[82] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[83] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[84] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[85] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[86] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[87] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[88] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[89] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[8] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[90] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[91] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[92] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[93] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[94] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[95] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[96] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[97] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[98] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[99] ;
 wire \Tile_X0Y1_DSP_bot/ConfigBits_N[9] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/E6BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/EE4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[0] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[10] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[11] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[12] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[13] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[14] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[15] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[16] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[17] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[18] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[19] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[1] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[20] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[21] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[22] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[23] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[24] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[25] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[26] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[27] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[28] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[29] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[2] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[30] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[31] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[3] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[4] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[5] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[6] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[7] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[8] ;
 wire \Tile_X0Y1_DSP_bot/FrameData_O_i[9] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[0] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[10] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[11] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[12] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[13] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[14] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[15] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[16] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[17] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[18] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[19] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[1] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[2] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[3] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[4] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[5] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[6] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[7] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[8] ;
 wire \Tile_X0Y1_DSP_bot/FrameStrobe_O_i[9] ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out2 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out3 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[0] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[10] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[11] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[12] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[13] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[14] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[15] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[16] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[17] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[18] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[19] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[1] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[2] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[3] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[4] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[5] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[6] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[7] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[8] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[9] ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0000_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0001_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0002_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0003_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0004_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0005_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0006_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0007_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0008_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0009_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0010_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0011_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0012_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0013_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0014_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0015_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0016_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0017_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0018_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0019_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0020_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0022_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0036_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0042_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0053_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0055_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0056_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0059_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0078_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0083_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0087_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0088_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0092_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0095_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0096_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0104_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0110_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0111_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0118_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0119_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0128_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0129_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0131_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0133_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0134_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0139_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0140_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0144_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0148_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0156_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0160_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0161_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0162_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0172_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0177_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0179_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0180_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0182_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0186_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0201_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0202_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0210_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0211_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0212_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0218_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0232_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0233_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0234_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0236_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0242_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0246_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0248_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0252_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0253_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0254_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0256_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0260_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0262_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0266_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0278_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0279_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0296_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0302_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0308_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0316_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0320_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0322_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0323_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0324_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0328_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0332_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0337_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0338_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0340_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0344_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0350_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0352_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0354_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0355_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0361_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0364_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0373_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0376_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0384_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0388_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0402_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0403_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0404_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0408_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0412_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0418_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0419_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0422_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0425_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0427_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0433_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0434_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0437_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0447_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0456_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0459_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0465_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0468_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0469_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0470_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0471_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0477_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0482_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0485_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0486_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0489_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0499_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0500_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0503_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0506_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0507_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0513_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0514_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0515_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0517_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0518_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0532_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0537_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0538_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0540_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0541_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0542_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0544_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0546_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0547_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0548_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0550_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0565_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0567_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0568_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0571_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0577_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0580_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0582_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0583_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0585_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0587_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0588_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0589_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0590_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0592_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0593_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0595_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0601_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0602_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0606_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0608_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0615_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0620_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0621_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0627_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0635_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0637_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0640_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0642_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0643_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0647_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0648_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0653_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0654_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0659_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0662_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0668_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0678_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0680_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0685_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0686_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0688_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0693_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0694_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0704_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0708_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0710_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0716_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0724_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0726_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0727_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0731_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0735_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0738_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0742_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0745_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0747_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0753_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0754_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0756_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0757_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0758_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0759_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0761_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0766_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0768_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0769_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0772_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0776_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0779_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0781_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0782_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0784_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0786_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0788_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0791_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0792_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0793_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0794_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0797_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0800_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0807_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0808_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0811_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0812_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0819_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0820_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0821_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0822_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0823_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0826_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0828_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0831_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0832_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0833_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0834_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0835_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0836_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0837_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0838_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0839_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0840_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0841_ ;
 wire \Tile_X0Y1_DSP_bot/Inst_MULADD/_0842_ ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JE2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JN2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JS2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[4] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[5] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[6] ;
 wire \Tile_X0Y1_DSP_bot/JW2BEG[7] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_AB_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_CD_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_EF_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[0] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[1] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[2] ;
 wire \Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/N4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/NN4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/Q0 ;
 wire \Tile_X0Y1_DSP_bot/Q1 ;
 wire \Tile_X0Y1_DSP_bot/Q10 ;
 wire \Tile_X0Y1_DSP_bot/Q11 ;
 wire \Tile_X0Y1_DSP_bot/Q12 ;
 wire \Tile_X0Y1_DSP_bot/Q13 ;
 wire \Tile_X0Y1_DSP_bot/Q14 ;
 wire \Tile_X0Y1_DSP_bot/Q15 ;
 wire \Tile_X0Y1_DSP_bot/Q16 ;
 wire \Tile_X0Y1_DSP_bot/Q17 ;
 wire \Tile_X0Y1_DSP_bot/Q18 ;
 wire \Tile_X0Y1_DSP_bot/Q19 ;
 wire \Tile_X0Y1_DSP_bot/Q2 ;
 wire \Tile_X0Y1_DSP_bot/Q3 ;
 wire \Tile_X0Y1_DSP_bot/Q4 ;
 wire \Tile_X0Y1_DSP_bot/Q5 ;
 wire \Tile_X0Y1_DSP_bot/Q6 ;
 wire \Tile_X0Y1_DSP_bot/Q7 ;
 wire \Tile_X0Y1_DSP_bot/Q8 ;
 wire \Tile_X0Y1_DSP_bot/Q9 ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/S4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/SS4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/W6BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[0] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[10] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[11] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[1] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[2] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[3] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[4] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[5] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[6] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[7] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[8] ;
 wire \Tile_X0Y1_DSP_bot/WW4BEG_i[9] ;
 wire \Tile_X0Y1_DSP_bot/clr ;
 wire \Tile_X0Y1_FrameStrobe_O[0] ;
 wire \Tile_X0Y1_FrameStrobe_O[10] ;
 wire \Tile_X0Y1_FrameStrobe_O[11] ;
 wire \Tile_X0Y1_FrameStrobe_O[12] ;
 wire \Tile_X0Y1_FrameStrobe_O[13] ;
 wire \Tile_X0Y1_FrameStrobe_O[14] ;
 wire \Tile_X0Y1_FrameStrobe_O[15] ;
 wire \Tile_X0Y1_FrameStrobe_O[16] ;
 wire \Tile_X0Y1_FrameStrobe_O[17] ;
 wire \Tile_X0Y1_FrameStrobe_O[18] ;
 wire \Tile_X0Y1_FrameStrobe_O[19] ;
 wire \Tile_X0Y1_FrameStrobe_O[1] ;
 wire \Tile_X0Y1_FrameStrobe_O[2] ;
 wire \Tile_X0Y1_FrameStrobe_O[3] ;
 wire \Tile_X0Y1_FrameStrobe_O[4] ;
 wire \Tile_X0Y1_FrameStrobe_O[5] ;
 wire \Tile_X0Y1_FrameStrobe_O[6] ;
 wire \Tile_X0Y1_FrameStrobe_O[7] ;
 wire \Tile_X0Y1_FrameStrobe_O[8] ;
 wire \Tile_X0Y1_FrameStrobe_O[9] ;
 wire \Tile_X0Y1_N1BEG[0] ;
 wire \Tile_X0Y1_N1BEG[1] ;
 wire \Tile_X0Y1_N1BEG[2] ;
 wire \Tile_X0Y1_N1BEG[3] ;
 wire \Tile_X0Y1_N2BEG[0] ;
 wire \Tile_X0Y1_N2BEG[1] ;
 wire \Tile_X0Y1_N2BEG[2] ;
 wire \Tile_X0Y1_N2BEG[3] ;
 wire \Tile_X0Y1_N2BEG[4] ;
 wire \Tile_X0Y1_N2BEG[5] ;
 wire \Tile_X0Y1_N2BEG[6] ;
 wire \Tile_X0Y1_N2BEG[7] ;
 wire \Tile_X0Y1_N2BEGb[0] ;
 wire \Tile_X0Y1_N2BEGb[1] ;
 wire \Tile_X0Y1_N2BEGb[2] ;
 wire \Tile_X0Y1_N2BEGb[3] ;
 wire \Tile_X0Y1_N2BEGb[4] ;
 wire \Tile_X0Y1_N2BEGb[5] ;
 wire \Tile_X0Y1_N2BEGb[6] ;
 wire \Tile_X0Y1_N2BEGb[7] ;
 wire \Tile_X0Y1_N4BEG[0] ;
 wire \Tile_X0Y1_N4BEG[10] ;
 wire \Tile_X0Y1_N4BEG[11] ;
 wire \Tile_X0Y1_N4BEG[12] ;
 wire \Tile_X0Y1_N4BEG[13] ;
 wire \Tile_X0Y1_N4BEG[14] ;
 wire \Tile_X0Y1_N4BEG[15] ;
 wire \Tile_X0Y1_N4BEG[1] ;
 wire \Tile_X0Y1_N4BEG[2] ;
 wire \Tile_X0Y1_N4BEG[3] ;
 wire \Tile_X0Y1_N4BEG[4] ;
 wire \Tile_X0Y1_N4BEG[5] ;
 wire \Tile_X0Y1_N4BEG[6] ;
 wire \Tile_X0Y1_N4BEG[7] ;
 wire \Tile_X0Y1_N4BEG[8] ;
 wire \Tile_X0Y1_N4BEG[9] ;
 wire \Tile_X0Y1_NN4BEG[0] ;
 wire \Tile_X0Y1_NN4BEG[10] ;
 wire \Tile_X0Y1_NN4BEG[11] ;
 wire \Tile_X0Y1_NN4BEG[12] ;
 wire \Tile_X0Y1_NN4BEG[13] ;
 wire \Tile_X0Y1_NN4BEG[14] ;
 wire \Tile_X0Y1_NN4BEG[15] ;
 wire \Tile_X0Y1_NN4BEG[1] ;
 wire \Tile_X0Y1_NN4BEG[2] ;
 wire \Tile_X0Y1_NN4BEG[3] ;
 wire \Tile_X0Y1_NN4BEG[4] ;
 wire \Tile_X0Y1_NN4BEG[5] ;
 wire \Tile_X0Y1_NN4BEG[6] ;
 wire \Tile_X0Y1_NN4BEG[7] ;
 wire \Tile_X0Y1_NN4BEG[8] ;
 wire \Tile_X0Y1_NN4BEG[9] ;
 wire Tile_X0Y1_UserCLKo;
 wire \Tile_X0Y1_bot2top[0] ;
 wire \Tile_X0Y1_bot2top[1] ;
 wire \Tile_X0Y1_bot2top[2] ;
 wire \Tile_X0Y1_bot2top[3] ;
 wire \Tile_X0Y1_bot2top[4] ;
 wire \Tile_X0Y1_bot2top[5] ;
 wire \Tile_X0Y1_bot2top[6] ;
 wire \Tile_X0Y1_bot2top[7] ;
 wire \Tile_X0Y1_bot2top[8] ;
 wire \Tile_X0Y1_bot2top[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\Tile_X0Y0_S1BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\Tile_X0Y0_SS4BEG[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\Tile_X0Y0_SS4BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\Tile_X0Y0_SS4BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\Tile_X0Y0_SS4BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(\Tile_X0Y0_SS4BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\Tile_X0Y1_FrameStrobe_O[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(\Tile_X0Y1_FrameStrobe_O[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\Tile_X0Y1_FrameStrobe_O[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\Tile_X0Y1_N1BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\Tile_X0Y0_DSP_top/E6BEG_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\Tile_X0Y0_DSP_top/SS4BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\Tile_X0Y0_DSP_top/SS4BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(\Tile_X0Y1_DSP_bot/E6BEG_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(\Tile_X0Y1_DSP_bot/N4BEG_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(\Tile_X0Y1_DSP_bot/S4BEG_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(\Tile_X0Y1_DSP_bot/SS4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\Tile_X0Y1_FrameStrobe_O[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\Tile_X0Y0_S1BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\Tile_X0Y1_FrameStrobe_O[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\Tile_X0Y0_S1BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\Tile_X0Y1_FrameStrobe_O[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\Tile_X0Y1_N1BEG[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\Tile_X0Y1_N2BEG[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\Tile_X0Y0_DSP_top/E6BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\Tile_X0Y0_DSP_top/EE4BEG_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\Tile_X0Y0_DSP_top/EE4BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\Tile_X0Y0_DSP_top/JE2BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\Tile_X0Y0_DSP_top/JE2BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\Tile_X0Y0_DSP_top/JN2BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\Tile_X0Y0_DSP_top/JS2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\Tile_X0Y0_SS4BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\Tile_X0Y0_DSP_top/JS2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\Tile_X0Y0_DSP_top/JS2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\Tile_X0Y0_DSP_top/JW2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\Tile_X0Y0_DSP_top/JW2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\Tile_X0Y0_DSP_top/JW2BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\Tile_X0Y0_DSP_top/JW2BEG[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\Tile_X0Y0_SS4BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\Tile_X0Y0_DSP_top/N4BEG_i[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\Tile_X0Y0_DSP_top/NN4BEG_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\Tile_X0Y0_SS4BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\Tile_X0Y0_DSP_top/S4BEG_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\Tile_X0Y0_DSP_top/W6BEG_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\Tile_X0Y1_DSP_bot/E6BEG_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\Tile_X0Y1_DSP_bot/EE4BEG_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\Tile_X0Y1_DSP_bot/JN2BEG[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\Tile_X0Y1_DSP_bot/N4BEG_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\Tile_X0Y1_DSP_bot/NN4BEG_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\Tile_X0Y1_DSP_bot/NN4BEG_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\Tile_X0Y1_DSP_bot/SS4BEG_i[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net144));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_91 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[0] ),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[1] ),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[2] ),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[3] ),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[4] ),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[5] ),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[6] ),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[7] ),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[8] ),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/E6BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/E6BEG_i[9] ),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_0/_0_  (.A(net25),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_1/_0_  (.A(net26),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_2/_0_  (.A(net27),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_3/_0_  (.A(net28),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_4/_0_  (.A(net29),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_5/_0_  (.A(net30),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_6/_0_  (.A(net31),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_7/_0_  (.A(net32),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_8/_0_  (.A(net22),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/E6END_inbuf_9/_0_  (.A(net23),
    .X(\Tile_X0Y0_DSP_top/E6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[0] ),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[1] ),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[10] ),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[11] ),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[2] ),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[3] ),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[4] ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[5] ),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[6] ),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[7] ),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[8] ),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/EE4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/EE4BEG_i[9] ),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_0/_0_  (.A(net43),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_1/_0_  (.A(net44),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_10/_0_  (.A(net38),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_11/_0_  (.A(net39),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_2/_0_  (.A(net45),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_3/_0_  (.A(net46),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_4/_0_  (.A(net47),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_5/_0_  (.A(net48),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_6/_0_  (.A(net34),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_7/_0_  (.A(net35),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_8/_0_  (.A(net36),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/EE4END_inbuf_9/_0_  (.A(net37),
    .X(\Tile_X0Y0_DSP_top/EE4BEG_i[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[374] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[375] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[384] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[385] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[386] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[387] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[388] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[389] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[390] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[391] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[392] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[393] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[376] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[394] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[395] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[396] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[397] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[398] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[399] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[400] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[401] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[402] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[403] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[377] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[404] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[405] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[378] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[378] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[379] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[380] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[381] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[382] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame0_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[0] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[383] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[54] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[55] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[64] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[65] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[66] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[67] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[68] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[69] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[70] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[71] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[72] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[73] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[56] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[74] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[75] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[76] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[77] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[78] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[79] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[80] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[81] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[82] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[83] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[57] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[84] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[85] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[58] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[59] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[60] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[61] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[62] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame10_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[10] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[63] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[22] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[23] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[32] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[33] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[34] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[35] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[36] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[37] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[38] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[39] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[40] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[41] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[24] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[42] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[43] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[44] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[45] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[46] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[47] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[50] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[51] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[25] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[26] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[27] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[28] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[29] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[30] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame11_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[11] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[31] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[0] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[1] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[2] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[3] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[4] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[5] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[6] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[7] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[8] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[9] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[10] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[11] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[12] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[13] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[14] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[15] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[16] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[17] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[18] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[19] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[20] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame12_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[12] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[21] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[352] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[353] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[356] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[357] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[360] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[361] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[344] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[364] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[365] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[368] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[369] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[345] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[372] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[373] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[348] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[349] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame1_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[1] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[320] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[321] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[324] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[325] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[328] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[329] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[312] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[332] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[333] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[336] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[337] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[313] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[340] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[341] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[316] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[317] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame2_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[2] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[288] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[289] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[292] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[293] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[296] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[297] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[280] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[300] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[301] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[304] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[305] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[281] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[308] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[309] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[284] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[285] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame3_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[3] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[256] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[257] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[260] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[261] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[264] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[265] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[248] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[268] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[269] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[272] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[273] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[249] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[276] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[277] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[252] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[253] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame4_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[4] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[214] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[215] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[224] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[225] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[226] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[227] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[228] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[229] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[230] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[231] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[232] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[233] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[216] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[234] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[235] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[236] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[237] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[238] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[239] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[240] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[241] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[242] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[243] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[217] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[244] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[245] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[218] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[219] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[220] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[221] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[222] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame5_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[5] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[223] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[182] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[183] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[192] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[193] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[194] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[195] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[196] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[197] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[198] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[199] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[200] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[201] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[184] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[202] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[203] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[204] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[205] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[206] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[207] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[208] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[209] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[210] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[211] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[185] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[212] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[213] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[186] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[187] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[188] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[189] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[190] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame6_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[6] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[191] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[150] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[151] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[160] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[161] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[162] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[163] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[164] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[165] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[166] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[167] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[168] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[169] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[152] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[170] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[171] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[172] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[173] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[174] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[175] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[176] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[177] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[178] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[179] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[153] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[180] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[181] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[154] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[155] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[156] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[157] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[158] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame7_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[7] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[159] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[118] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[119] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[128] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[129] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[130] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[131] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[132] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[133] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[134] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[135] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[136] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[137] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[120] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[138] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[139] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[140] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[141] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[142] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[143] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[144] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[145] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[146] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[147] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[121] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[148] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[149] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[122] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[123] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[124] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[125] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[126] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame8_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[8] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[127] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit0  (.D(net49),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[86] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit1  (.D(net60),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[87] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit10  (.D(net50),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[96] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit11  (.D(net51),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[97] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit12  (.D(net52),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[98] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit13  (.D(net53),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[99] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit14  (.D(net54),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[100] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit15  (.D(net55),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[101] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit16  (.D(net56),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[102] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit17  (.D(net57),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[103] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit18  (.D(net58),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit19  (.D(net59),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit2  (.D(net71),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[88] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit20  (.D(net61),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[106] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit21  (.D(net62),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[107] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit22  (.D(net63),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit23  (.D(net64),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit24  (.D(net65),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[110] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit25  (.D(net66),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[111] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit26  (.D(net67),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[112] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit27  (.D(net68),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[113] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit28  (.D(net69),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[114] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit29  (.D(net70),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[115] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit3  (.D(net74),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[89] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit30  (.D(net72),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[116] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit31  (.D(net73),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[117] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit4  (.D(net75),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[90] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit5  (.D(net76),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[91] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit6  (.D(net77),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[92] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit7  (.D(net78),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[93] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit8  (.D(net79),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[94] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_ConfigMem/Inst_frame9_bit9  (.D(net80),
    .GATE(\Tile_X0Y1_FrameStrobe_O[9] ),
    .Q(\Tile_X0Y0_DSP_top/ConfigBits[95] ),
    .Q_N(\Tile_X0Y0_DSP_top/ConfigBits_N[95] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_00_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[0] ),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_01_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[1] ),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_02_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[2] ),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_03_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_04_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_05_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[5] ),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_06_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[6] ),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_07_  (.A(\Tile_X0Y0_DSP_top/JE2BEG[7] ),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_08_  (.A(net13),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_09_  (.A(net14),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_10_  (.A(net15),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_11_  (.A(net16),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_12_  (.A(net17),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_13_  (.A(net18),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_14_  (.A(net19),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_15_  (.A(net20),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_16_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[0] ),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_17_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[1] ),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_18_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_19_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_20_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_21_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[5] ),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_22_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[6] ),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_23_  (.A(\Tile_X0Y0_DSP_top/JN2BEG[7] ),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_24_  (.A(\Tile_X0Y1_N2BEG[0] ),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_25_  (.A(\Tile_X0Y1_N2BEG[1] ),
    .X(net495));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_26_  (.A(\Tile_X0Y1_N2BEG[2] ),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_27_  (.A(\Tile_X0Y1_N2BEG[3] ),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_28_  (.A(\Tile_X0Y1_N2BEG[4] ),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_29_  (.A(\Tile_X0Y1_N2BEG[5] ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_30_  (.A(\Tile_X0Y1_N2BEG[6] ),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_31_  (.A(\Tile_X0Y1_N2BEG[7] ),
    .X(net501));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_32_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[0] ),
    .X(\Tile_X0Y0_S2BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_33_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[1] ),
    .X(\Tile_X0Y0_S2BEG[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_34_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[2] ),
    .X(\Tile_X0Y0_S2BEG[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_35_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .X(\Tile_X0Y0_S2BEG[3] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_36_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .X(\Tile_X0Y0_S2BEG[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_37_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[5] ),
    .X(\Tile_X0Y0_S2BEG[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_38_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[6] ),
    .X(\Tile_X0Y0_S2BEG[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_39_  (.A(\Tile_X0Y0_DSP_top/JS2BEG[7] ),
    .X(\Tile_X0Y0_S2BEG[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_40_  (.A(net93),
    .X(\Tile_X0Y0_S2BEGb[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_41_  (.A(net94),
    .X(\Tile_X0Y0_S2BEGb[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_42_  (.A(net95),
    .X(\Tile_X0Y0_S2BEGb[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_43_  (.A(net96),
    .X(\Tile_X0Y0_S2BEGb[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_44_  (.A(net97),
    .X(\Tile_X0Y0_S2BEGb[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_45_  (.A(net98),
    .X(\Tile_X0Y0_S2BEGb[5] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_46_  (.A(net99),
    .X(\Tile_X0Y0_S2BEGb[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_47_  (.A(net100),
    .X(\Tile_X0Y0_S2BEGb[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_48_  (.A(net137),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_49_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[1] ),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_50_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[2] ),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_51_  (.A(net140),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_52_  (.A(net141),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_53_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[5] ),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_54_  (.A(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_55_  (.A(net144),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_56_  (.A(net145),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_57_  (.A(net146),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_58_  (.A(net147),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_59_  (.A(net148),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_60_  (.A(net149),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_61_  (.A(net150),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_62_  (.A(net151),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/_63_  (.A(net152),
    .X(net554));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net136),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[48] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[49] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[50] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[51] ),
    .X(net403));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0  (.A0(net3),
    .A1(net135),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[52] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[53] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[54] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[55] ),
    .X(net404));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[1] ),
    .A2(\Tile_X0Y1_N4BEG[1] ),
    .A3(net40),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net86),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[278] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[279] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[280] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[281] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[2] ),
    .A2(\Tile_X0Y1_N4BEG[2] ),
    .A3(net7),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net87),
    .A2(net139),
    .A3(net174),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[282] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[283] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[284] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[285] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[3] ),
    .A2(\Tile_X0Y1_N4BEG[3] ),
    .A3(net8),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net88),
    .A2(net140),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[286] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[287] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[288] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[289] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[4] ),
    .A2(\Tile_X0Y1_N4BEG[0] ),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net89),
    .A2(net141),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[290] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[291] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[292] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[293] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net90),
    .A3(net134),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[294] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[295] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[296] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[297] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net91),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[298] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[299] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[300] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[301] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net92),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[302] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[303] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[304] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[305] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net117),
    .A3(net165),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[306] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[307] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[308] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[309] ),
    .X(\Tile_X0Y0_DSP_top/JE2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[1] ),
    .A1(\Tile_X0Y1_N4BEG[1] ),
    .A2(net4),
    .A3(net6),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net124),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[246] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[247] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[248] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[249] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[2] ),
    .A1(\Tile_X0Y1_N4BEG[2] ),
    .A2(net1),
    .A3(net7),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net87),
    .A2(net139),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[250] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[251] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[252] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[253] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(\Tile_X0Y1_N4BEG[3] ),
    .A2(net2),
    .A3(net8),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1  (.A0(net24),
    .A1(net88),
    .A2(net140),
    .A3(net172),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[254] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[255] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[256] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[257] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(\Tile_X0Y1_N4BEG[0] ),
    .A2(net3),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1  (.A0(net21),
    .A1(net89),
    .A2(net141),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[258] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[259] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[260] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[261] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net90),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[262] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[263] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[264] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[265] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1  (.A0(net83),
    .A1(net91),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[266] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[267] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[268] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[269] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1  (.A0(net84),
    .A1(net92),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[270] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[271] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[272] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[273] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net33),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net85),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[274] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[275] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[276] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[277] ),
    .X(\Tile_X0Y0_DSP_top/JN2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_NN4BEG[1] ),
    .A1(net4),
    .A2(net6),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1  (.A0(net86),
    .A1(net108),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[310] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[311] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[312] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[313] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_NN4BEG[2] ),
    .A1(net1),
    .A2(net41),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1  (.A0(net109),
    .A1(net125),
    .A2(net139),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[314] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[315] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[316] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[317] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_NN4BEG[3] ),
    .A1(net2),
    .A2(net8),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1  (.A0(net88),
    .A1(net110),
    .A2(net140),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[318] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[319] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[320] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[321] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(net3),
    .A2(net9),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1  (.A0(net89),
    .A1(net101),
    .A2(net141),
    .A3(net173),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[322] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[323] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[324] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[325] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net90),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[326] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[327] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[328] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[329] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1  (.A0(net83),
    .A1(net91),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[330] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[331] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[332] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[333] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1  (.A0(net84),
    .A1(net92),
    .A2(net134),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[334] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[335] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[336] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[337] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net85),
    .A2(net133),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[338] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[339] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[340] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[341] ),
    .X(\Tile_X0Y0_DSP_top/JS2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[1] ),
    .A2(net6),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1  (.A0(net86),
    .A1(net108),
    .A2(net138),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[1] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[342] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[343] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[344] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[345] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[2] ),
    .A2(net7),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1  (.A0(net87),
    .A1(net109),
    .A2(net139),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[2] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[346] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[347] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[348] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[349] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[3] ),
    .A2(net8),
    .A3(net24),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1  (.A0(net88),
    .A1(net110),
    .A2(net140),
    .A3(net156),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[3] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[350] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[351] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[352] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[353] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[4] ),
    .A2(net9),
    .A3(net21),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1  (.A0(net89),
    .A1(net101),
    .A2(net141),
    .A3(net153),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[354] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[355] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[356] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[357] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(\Tile_X0Y1_N2BEGb[5] ),
    .A2(net2),
    .A3(net10),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net90),
    .A3(net134),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[358] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[359] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[360] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[361] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(\Tile_X0Y1_N2BEGb[6] ),
    .A2(net3),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net91),
    .A3(net135),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[6] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[362] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[363] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[364] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[365] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(\Tile_X0Y1_N2BEGb[7] ),
    .A2(net4),
    .A3(net12),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1  (.A0(net82),
    .A1(net84),
    .A2(net92),
    .A3(net136),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[7] ),
    .A3(\Tile_X0Y1_bot2top[8] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[366] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[367] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[368] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[369] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(\Tile_X0Y1_N2BEGb[0] ),
    .A2(net1),
    .A3(net5),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1  (.A0(net81),
    .A1(net83),
    .A2(net85),
    .A3(net133),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y1_bot2top[1] ),
    .A2(\Tile_X0Y1_bot2top[2] ),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y1_bot2top[5] ),
    .A2(\Tile_X0Y1_bot2top[6] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[370] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[371] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[372] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[373] ),
    .X(\Tile_X0Y0_DSP_top/JW2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net136),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[104] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[105] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[106] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[107] ),
    .X(net556));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0  (.A0(net3),
    .A1(net135),
    .A2(\Tile_X0Y1_bot2top[0] ),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y1_bot2top[3] ),
    .A2(\Tile_X0Y1_bot2top[4] ),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y1_bot2top[7] ),
    .A2(\Tile_X0Y1_bot2top[8] ),
    .A3(\Tile_X0Y1_bot2top[9] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[108] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[109] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[110] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[111] ),
    .X(net557));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG0  (.A0(\Tile_X0Y1_bot2top[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[28] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[29] ),
    .X(net382));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG1  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[30] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[31] ),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG2  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[32] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[33] ),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_E1BEG3  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[34] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[35] ),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(\Tile_X0Y1_N2BEGb[6] ),
    .A1(net11),
    .A2(net126),
    .A3(net143),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[214] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[215] ),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(\Tile_X0Y1_NN4BEG[0] ),
    .A1(net7),
    .A2(net87),
    .A3(net139),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[216] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[217] ),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(net33),
    .A2(net89),
    .A3(net141),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[218] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[219] ),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(\Tile_X0Y1_N2BEGb[0] ),
    .A1(net5),
    .A2(net85),
    .A3(net174),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[220] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[221] ),
    .X(\Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(\Tile_X0Y1_NN4BEG[3] ),
    .A1(net11),
    .A2(net91),
    .A3(net143),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[222] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[223] ),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(\Tile_X0Y1_N2BEGb[2] ),
    .A1(net7),
    .A2(net87),
    .A3(net173),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[224] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[225] ),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(\Tile_X0Y1_N2BEGb[4] ),
    .A1(net9),
    .A2(net125),
    .A3(net141),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[226] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[227] ),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(\Tile_X0Y1_N2BEGb[0] ),
    .A1(net40),
    .A2(net85),
    .A3(net137),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[228] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[229] ),
    .X(\Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(\Tile_X0Y1_N2BEGb[7] ),
    .A1(net41),
    .A2(net92),
    .A3(net144),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[230] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[231] ),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(net8),
    .A2(net88),
    .A3(net172),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[232] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[233] ),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(\Tile_X0Y1_N2BEGb[5] ),
    .A1(net10),
    .A2(net124),
    .A3(net142),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[234] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[235] ),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(\Tile_X0Y1_NN4BEG[2] ),
    .A1(net6),
    .A2(net86),
    .A3(net138),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[236] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[237] ),
    .X(\Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(\Tile_X0Y1_N2BEGb[7] ),
    .A1(net12),
    .A2(net92),
    .A3(net165),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[238] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[239] ),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(net8),
    .A2(net117),
    .A3(net140),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[240] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[241] ),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(\Tile_X0Y1_NN4BEG[1] ),
    .A1(net10),
    .A2(net90),
    .A3(net142),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[242] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[243] ),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(\Tile_X0Y1_N2BEGb[1] ),
    .A1(net42),
    .A2(net86),
    .A3(net138),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[244] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[245] ),
    .X(\Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(\Tile_X0Y1_N2BEG[6] ),
    .A1(net99),
    .A2(net151),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[150] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[151] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net15),
    .A1(net95),
    .A2(net147),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[152] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[153] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(\Tile_X0Y1_N2BEG[4] ),
    .A1(net17),
    .A2(net149),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[154] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[155] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(\Tile_X0Y1_N2BEG[0] ),
    .A1(net13),
    .A2(net93),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[156] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[157] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[182] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[183] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[184] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[185] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[186] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[187] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[188] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[189] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net19),
    .A1(net99),
    .A2(net151),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[158] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[159] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(\Tile_X0Y1_N2BEG[2] ),
    .A1(net15),
    .A2(net147),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[160] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[161] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(\Tile_X0Y1_N2BEG[4] ),
    .A1(net17),
    .A2(net97),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[162] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[163] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(\Tile_X0Y1_N2BEG[0] ),
    .A1(net93),
    .A2(net145),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[164] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[165] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[190] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[191] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[192] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[193] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[194] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[195] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[196] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[197] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(\Tile_X0Y1_N2BEG[6] ),
    .A1(net19),
    .A2(net151),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[166] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[167] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(\Tile_X0Y1_N2BEG[2] ),
    .A1(net15),
    .A2(net95),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[168] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[169] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(\Tile_X0Y1_N2BEG[4] ),
    .A1(net97),
    .A2(net149),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[170] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[171] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net13),
    .A1(net93),
    .A2(net145),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[172] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[173] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[198] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[199] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[200] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[201] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[202] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[203] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[204] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[205] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(\Tile_X0Y1_N2BEG[6] ),
    .A1(net19),
    .A2(net99),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[174] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[175] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(\Tile_X0Y1_N2BEG[2] ),
    .A1(net95),
    .A2(net147),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[176] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[177] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net17),
    .A1(net97),
    .A2(net149),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[178] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[179] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(\Tile_X0Y1_N2BEG[0] ),
    .A1(net13),
    .A2(net145),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[180] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[181] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(\Tile_X0Y1_N2BEG[7] ),
    .A1(net20),
    .A2(net100),
    .A3(net152),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[206] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[207] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(\Tile_X0Y1_N2BEG[3] ),
    .A1(net16),
    .A2(net96),
    .A3(net148),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[208] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[209] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(\Tile_X0Y1_N2BEG[5] ),
    .A1(net18),
    .A2(net98),
    .A3(net150),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[210] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[211] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(\Tile_X0Y1_N2BEG[1] ),
    .A1(net14),
    .A2(net94),
    .A3(net146),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[212] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[213] ),
    .X(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(\Tile_X0Y1_NN4BEG[3] ),
    .A1(net110),
    .A2(net165),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[374] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[375] ),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net41),
    .A1(net109),
    .A2(net144),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[376] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[377] ),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(\Tile_X0Y1_N4BEG[1] ),
    .A1(net24),
    .A2(net156),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[378] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[379] ),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(\Tile_X0Y1_N4BEG[0] ),
    .A1(net21),
    .A2(net101),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[380] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[381] ),
    .X(\Tile_X0Y0_DSP_top/J_l_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net8),
    .A1(net126),
    .A2(net173),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[382] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[383] ),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(\Tile_X0Y1_N4BEG[2] ),
    .A1(net7),
    .A2(net144),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[384] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[385] ),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(\Tile_X0Y1_NN4BEG[1] ),
    .A1(net40),
    .A2(net108),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[386] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[387] ),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(\Tile_X0Y1_N4BEG[0] ),
    .A1(net117),
    .A2(net153),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[388] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[389] ),
    .X(\Tile_X0Y0_DSP_top/J_l_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(\Tile_X0Y1_N4BEG[3] ),
    .A1(net8),
    .A2(net140),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[390] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[391] ),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(\Tile_X0Y1_NN4BEG[2] ),
    .A1(net7),
    .A2(net109),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[392] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[393] ),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(\Tile_X0Y1_N4BEG[1] ),
    .A1(net124),
    .A2(net141),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[394] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[395] ),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net42),
    .A1(net101),
    .A2(net172),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[396] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[397] ),
    .X(\Tile_X0Y0_DSP_top/J_l_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(\Tile_X0Y1_N4BEG[3] ),
    .A1(net33),
    .A2(net110),
    .A3(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[398] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[399] ),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(\Tile_X0Y1_N4BEG[2] ),
    .A1(net125),
    .A2(net139),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[400] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[401] ),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net24),
    .A1(net108),
    .A2(net174),
    .A3(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[402] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[403] ),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(\Tile_X0Y1_NN4BEG[0] ),
    .A1(net21),
    .A2(net137),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[404] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[405] ),
    .X(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(\Tile_X0Y1_bot2top[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[0] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[1] ),
    .X(net482));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(\Tile_X0Y1_bot2top[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[2] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[3] ),
    .X(net483));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[4] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[5] ),
    .X(net484));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[6] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[7] ),
    .X(net485));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG0  (.A0(\Tile_X0Y1_N2BEGb[2] ),
    .A1(\Tile_X0Y1_N4BEG[1] ),
    .A2(net24),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[8] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[9] ),
    .X(net505));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG1  (.A0(\Tile_X0Y1_N2BEGb[3] ),
    .A1(\Tile_X0Y1_N4BEG[2] ),
    .A2(net21),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[10] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[11] ),
    .X(net506));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG2  (.A0(\Tile_X0Y1_N2BEGb[0] ),
    .A1(\Tile_X0Y1_N4BEG[3] ),
    .A2(net156),
    .A3(\Tile_X0Y1_bot2top[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[12] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[13] ),
    .X(net507));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_N4BEG3  (.A0(\Tile_X0Y1_N2BEGb[1] ),
    .A1(\Tile_X0Y1_N4BEG[0] ),
    .A2(net153),
    .A3(\Tile_X0Y1_bot2top[7] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[14] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[15] ),
    .X(net508));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(\Tile_X0Y1_bot2top[4] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[56] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[57] ),
    .X(\Tile_X0Y0_S1BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[58] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[59] ),
    .X(\Tile_X0Y0_S1BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[60] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[61] ),
    .X(\Tile_X0Y0_S1BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[62] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[63] ),
    .X(\Tile_X0Y0_S1BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG0  (.A0(net24),
    .A1(net87),
    .A2(net108),
    .A3(\Tile_X0Y1_bot2top[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[64] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[65] ),
    .X(\Tile_X0Y0_S4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG1  (.A0(net21),
    .A1(net88),
    .A2(net109),
    .A3(\Tile_X0Y1_bot2top[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[66] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[67] ),
    .X(\Tile_X0Y0_S4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG2  (.A0(net85),
    .A1(net110),
    .A2(net156),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[68] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[69] ),
    .X(\Tile_X0Y0_S4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_S4BEG3  (.A0(net86),
    .A1(net101),
    .A2(net153),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[70] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[71] ),
    .X(\Tile_X0Y0_S4BEG[15] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(\Tile_X0Y1_bot2top[5] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[84] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[85] ),
    .X(net535));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[86] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[87] ),
    .X(net536));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[88] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[89] ),
    .X(net537));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(\Tile_X0Y1_bot2top[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/JS2BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[90] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[91] ),
    .X(net538));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot0  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[112] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[113] ),
    .X(\Tile_X0Y0_top2bot[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot1  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[114] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[115] ),
    .X(\Tile_X0Y0_top2bot[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot10  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[132] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[133] ),
    .X(\Tile_X0Y0_top2bot[10] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot11  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[134] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[135] ),
    .X(\Tile_X0Y0_top2bot[11] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot12  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[136] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[137] ),
    .X(\Tile_X0Y0_top2bot[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot13  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[138] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[139] ),
    .X(\Tile_X0Y0_top2bot[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot14  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[140] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[141] ),
    .X(\Tile_X0Y0_top2bot[14] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot15  (.A0(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[142] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[143] ),
    .X(\Tile_X0Y0_top2bot[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot2  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[116] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[117] ),
    .X(\Tile_X0Y0_top2bot[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot3  (.A0(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_AB_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[118] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[119] ),
    .X(\Tile_X0Y0_top2bot[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot4  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[120] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[121] ),
    .X(\Tile_X0Y0_top2bot[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot5  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[122] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[123] ),
    .X(\Tile_X0Y0_top2bot[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot6  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[124] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[125] ),
    .X(\Tile_X0Y0_top2bot[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot7  (.A0(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[3] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_CD_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[126] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[127] ),
    .X(\Tile_X0Y0_top2bot[7] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot8  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[0] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[128] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[129] ),
    .X(\Tile_X0Y0_top2bot[8] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux41_buf_top2bot9  (.A0(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[1] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J_l_EF_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[130] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[131] ),
    .X(\Tile_X0Y0_top2bot[9] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net3),
    .A2(net83),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[36] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[37] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[36] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[37] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[38] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[38] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ),
    .Y(net417));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net4),
    .A2(net84),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[39] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[40] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[39] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[40] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[41] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[41] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ),
    .Y(net418));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net1),
    .A2(net81),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[42] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[43] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[42] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[43] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[44] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[44] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ),
    .Y(net419));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net2),
    .A2(net82),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[45] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[46] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[0] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[45] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[46] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[47] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[47] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ),
    .Y(net420));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net3),
    .A2(net135),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[16] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[17] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[16] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[17] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[18] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[18] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ),
    .Y(net521));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net4),
    .A2(net136),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[19] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[20] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[19] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[20] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[21] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[21] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ),
    .Y(net522));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net1),
    .A2(net133),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[22] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[23] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[22] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[23] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[24] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[24] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ),
    .Y(net523));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net2),
    .A2(net134),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[25] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[26] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[1] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[25] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[26] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[27] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[27] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ),
    .Y(net524));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net3),
    .A2(net135),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[72] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[73] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[72] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[73] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[74] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[74] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y0_SS4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net4),
    .A2(net136),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[75] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[76] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[75] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[76] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[77] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[77] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y0_SS4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net1),
    .A2(net133),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[78] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[79] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[78] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[79] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[80] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[80] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y0_SS4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net2),
    .A2(net134),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[81] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[82] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[81] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[82] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[83] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[83] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y0_SS4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[2] ),
    .A1(net83),
    .A2(net135),
    .A3(\Tile_X0Y1_bot2top[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[92] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[93] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[6] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_GH_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[92] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[93] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[94] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[94] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ),
    .Y(net570));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[3] ),
    .A1(net84),
    .A2(net136),
    .A3(\Tile_X0Y1_bot2top[3] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[95] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[96] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[7] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_EF_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[95] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[96] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[97] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[97] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ),
    .Y(net571));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[0] ),
    .A1(net81),
    .A2(net133),
    .A3(\Tile_X0Y1_bot2top[4] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[98] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[99] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[8] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_CD_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[98] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[99] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[100] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[100] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ),
    .Y(net572));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_N1BEG[1] ),
    .A1(net82),
    .A2(net134),
    .A3(\Tile_X0Y1_bot2top[5] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[101] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[102] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_bot2top[9] ),
    .A1(\Tile_X0Y0_DSP_top/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y0_DSP_top/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y0_DSP_top/J2END_AB_BEG[2] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[101] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[102] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[103] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[103] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ),
    .Y(net573));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_inst0  (.A0(\Tile_X0Y0_DSP_top/JN2BEG[4] ),
    .A1(\Tile_X0Y0_DSP_top/JN2BEG[6] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[4] ),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[144] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[145] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_DSP_top/JS2BEG[4] ),
    .A1(\Tile_X0Y0_DSP_top/JS2BEG[6] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[4] ),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[6] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[144] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[145] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[146] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[146] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot16/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y0_top2bot[16] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_inst0  (.A0(\Tile_X0Y0_DSP_top/JN2BEG[5] ),
    .A1(\Tile_X0Y0_DSP_top/JN2BEG[7] ),
    .A2(\Tile_X0Y0_DSP_top/JE2BEG[5] ),
    .A3(\Tile_X0Y0_DSP_top/JE2BEG[7] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[147] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[148] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_DSP_top/JS2BEG[5] ),
    .A1(\Tile_X0Y0_DSP_top/JS2BEG[7] ),
    .A2(\Tile_X0Y0_DSP_top/JW2BEG[5] ),
    .A3(\Tile_X0Y0_DSP_top/JW2BEG[7] ),
    .S0(\Tile_X0Y0_DSP_top/ConfigBits[147] ),
    .S1(\Tile_X0Y0_DSP_top/ConfigBits[148] ),
    .X(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_2_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_3_  (.A(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y0_DSP_top/ConfigBits[149] ),
    .Y(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_4_  (.A1(\Tile_X0Y0_DSP_top/ConfigBits[149] ),
    .A2(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y0_DSP_top/Inst_DSP_top_switch_matrix/inst_cus_mux81_buf_top2bot17/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y0_top2bot[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[0] ),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[1] ),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[10] ),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[11] ),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[2] ),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[3] ),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[4] ),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[5] ),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[6] ),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[7] ),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[8] ),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/N4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/N4BEG_i[9] ),
    .X(net517));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_0/_0_  (.A(\Tile_X0Y1_N4BEG[4] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_1/_0_  (.A(\Tile_X0Y1_N4BEG[5] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/N4END_inbuf_10/_0_  (.A(\Tile_X0Y1_N4BEG[14] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/N4END_inbuf_11/_0_  (.A(\Tile_X0Y1_N4BEG[15] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_2/_0_  (.A(\Tile_X0Y1_N4BEG[6] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_3/_0_  (.A(\Tile_X0Y1_N4BEG[7] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[3] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_4/_0_  (.A(\Tile_X0Y1_N4BEG[8] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[4] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_5/_0_  (.A(\Tile_X0Y1_N4BEG[9] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[5] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_6/_0_  (.A(\Tile_X0Y1_N4BEG[10] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_7/_0_  (.A(\Tile_X0Y1_N4BEG[11] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/N4END_inbuf_8/_0_  (.A(\Tile_X0Y1_N4BEG[12] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[8] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/N4END_inbuf_9/_0_  (.A(\Tile_X0Y1_N4BEG[13] ),
    .X(\Tile_X0Y0_DSP_top/N4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[0] ),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[1] ),
    .X(net525));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[10] ),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[11] ),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[2] ),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[3] ),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[4] ),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[5] ),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[6] ),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[7] ),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[8] ),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/NN4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/NN4BEG_i[9] ),
    .X(net533));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_0/_0_  (.A(\Tile_X0Y1_NN4BEG[4] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_1/_0_  (.A(\Tile_X0Y1_NN4BEG[5] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_10/_0_  (.A(\Tile_X0Y1_NN4BEG[14] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[10] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_11/_0_  (.A(\Tile_X0Y1_NN4BEG[15] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_2/_0_  (.A(\Tile_X0Y1_NN4BEG[6] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_3/_0_  (.A(\Tile_X0Y1_NN4BEG[7] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_4/_0_  (.A(\Tile_X0Y1_NN4BEG[8] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[4] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_5/_0_  (.A(\Tile_X0Y1_NN4BEG[9] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_6/_0_  (.A(\Tile_X0Y1_NN4BEG[10] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_7/_0_  (.A(\Tile_X0Y1_NN4BEG[11] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/NN4END_inbuf_8/_0_  (.A(\Tile_X0Y1_NN4BEG[12] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/NN4END_inbuf_9/_0_  (.A(\Tile_X0Y1_NN4BEG[13] ),
    .X(\Tile_X0Y0_DSP_top/NN4BEG_i[9] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[0] ),
    .X(\Tile_X0Y0_S4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[1] ),
    .X(\Tile_X0Y0_S4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[10] ),
    .X(\Tile_X0Y0_S4BEG[10] ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y0_DSP_top/S4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[11] ),
    .X(\Tile_X0Y0_S4BEG[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[2] ),
    .X(\Tile_X0Y0_S4BEG[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[3] ),
    .X(\Tile_X0Y0_S4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[4] ),
    .X(\Tile_X0Y0_S4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[5] ),
    .X(\Tile_X0Y0_S4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[6] ),
    .X(\Tile_X0Y0_S4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[7] ),
    .X(\Tile_X0Y0_S4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[8] ),
    .X(\Tile_X0Y0_S4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/S4BEG_i[9] ),
    .X(\Tile_X0Y0_S4BEG[9] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_0/_0_  (.A(net111),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_1/_0_  (.A(net112),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_10/_0_  (.A(net106),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/S4END_inbuf_11/_0_  (.A(net107),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_2/_0_  (.A(net113),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_3/_0_  (.A(net114),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_4/_0_  (.A(net115),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_5/_0_  (.A(net116),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_6/_0_  (.A(net102),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_7/_0_  (.A(net103),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/S4END_inbuf_8/_0_  (.A(net104),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/S4END_inbuf_9/_0_  (.A(net105),
    .X(\Tile_X0Y0_DSP_top/S4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[0] ),
    .X(\Tile_X0Y0_SS4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[1] ),
    .X(\Tile_X0Y0_SS4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[10] ),
    .X(\Tile_X0Y0_SS4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[11] ),
    .X(\Tile_X0Y0_SS4BEG[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[2] ),
    .X(\Tile_X0Y0_SS4BEG[2] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[3] ),
    .X(\Tile_X0Y0_SS4BEG[3] ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[4] ),
    .X(\Tile_X0Y0_SS4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[5] ),
    .X(\Tile_X0Y0_SS4BEG[5] ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[6] ),
    .X(\Tile_X0Y0_SS4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[7] ),
    .X(\Tile_X0Y0_SS4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[8] ),
    .X(\Tile_X0Y0_SS4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/SS4BEG_i[9] ),
    .X(\Tile_X0Y0_SS4BEG[9] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4END_inbuf_0/_0_  (.A(net127),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y0_DSP_top/SS4END_inbuf_1/_0_  (.A(net128),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_10/_0_  (.A(net122),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_11/_0_  (.A(net123),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y0_DSP_top/SS4END_inbuf_2/_0_  (.A(net129),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_3/_0_  (.A(net130),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_4/_0_  (.A(net131),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_5/_0_  (.A(net132),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_6/_0_  (.A(net118),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_7/_0_  (.A(net119),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_8/_0_  (.A(net120),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/SS4END_inbuf_9/_0_  (.A(net121),
    .X(\Tile_X0Y0_DSP_top/SS4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[0] ),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[1] ),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[2] ),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[3] ),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[4] ),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[5] ),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[6] ),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[7] ),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[8] ),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/W6BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/W6BEG_i[9] ),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_0/_0_  (.A(net157),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_1/_0_  (.A(net158),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_2/_0_  (.A(net159),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_3/_0_  (.A(net160),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_4/_0_  (.A(net161),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_5/_0_  (.A(net162),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_6/_0_  (.A(net163),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_7/_0_  (.A(net164),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_8/_0_  (.A(net154),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/W6END_inbuf_9/_0_  (.A(net155),
    .X(\Tile_X0Y0_DSP_top/W6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[0] ),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[1] ),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[10] ),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[11] ),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[2] ),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[3] ),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[4] ),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[5] ),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[6] ),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[7] ),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[8] ),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/WW4BEG_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/WW4BEG_i[9] ),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_0/_0_  (.A(net175),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_1/_0_  (.A(net176),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_10/_0_  (.A(net170),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_11/_0_  (.A(net171),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_2/_0_  (.A(net177),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_3/_0_  (.A(net178),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_4/_0_  (.A(net179),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_5/_0_  (.A(net180),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_6/_0_  (.A(net166),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_7/_0_  (.A(net167),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_8/_0_  (.A(net168),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y0_DSP_top/WW4END_inbuf_9/_0_  (.A(net169),
    .X(\Tile_X0Y0_DSP_top/WW4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_0/_0_  (.A(net49),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_1/_0_  (.A(net60),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_10/_0_  (.A(net50),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_11/_0_  (.A(net51),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_12/_0_  (.A(net52),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_13/_0_  (.A(net53),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_14/_0_  (.A(net54),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_15/_0_  (.A(net55),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_16/_0_  (.A(net56),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[16] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_17/_0_  (.A(net57),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_18/_0_  (.A(net58),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_19/_0_  (.A(net59),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_2/_0_  (.A(net71),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_20/_0_  (.A(net61),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[20] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_21/_0_  (.A(net62),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_22/_0_  (.A(net63),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_23/_0_  (.A(net64),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_24/_0_  (.A(net65),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_25/_0_  (.A(net66),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_26/_0_  (.A(net67),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_27/_0_  (.A(net68),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_28/_0_  (.A(net69),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_29/_0_  (.A(net70),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_3/_0_  (.A(net74),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[3] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_30/_0_  (.A(net72),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[30] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_inbuf_31/_0_  (.A(net73),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_4/_0_  (.A(net75),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_5/_0_  (.A(net76),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_6/_0_  (.A(net77),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_7/_0_  (.A(net78),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_8/_0_  (.A(net79),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_inbuf_9/_0_  (.A(net80),
    .X(\Tile_X0Y0_DSP_top/FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[0] ),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[1] ),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[10] ),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[11] ),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_12/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[12] ),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_13/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[13] ),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_14/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[14] ),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_15/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[15] ),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_16/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[16] ),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_17/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[17] ),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_18/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[18] ),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_19/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[19] ),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[2] ),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_20/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[20] ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_21/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[21] ),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_22/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[22] ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_23/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[23] ),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_24/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[24] ),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_25/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[25] ),
    .X(net447));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/data_outbuf_26/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[26] ),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_27/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[27] ),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_28/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[28] ),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_29/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[29] ),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[3] ),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_30/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[30] ),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_31/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[31] ),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[4] ),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[5] ),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[6] ),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[7] ),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[8] ),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/data_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/FrameData_O_i[9] ),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/inst_clk_buf  (.A(Tile_X0Y1_UserCLKo),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_0/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[0] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_1/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[1] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_10/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[10] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_11/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[11] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_12/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[12] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_13/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[13] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_14/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[14] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_15/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[15] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_16/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[16] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_17/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[17] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_18/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[18] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_19/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[19] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_2/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[2] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_3/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[3] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_4/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[4] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_5/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[5] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_6/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[6] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_7/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[7] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_8/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[8] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_inbuf_9/_0_  (.A(\Tile_X0Y1_FrameStrobe_O[9] ),
    .X(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_0/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[0] ),
    .X(net462));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_1/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[1] ),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_10/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[10] ),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_11/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[11] ),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_12/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[12] ),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_13/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[13] ),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_14/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[14] ),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_15/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[15] ),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_16/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[16] ),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_17/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[17] ),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_18/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[18] ),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_19/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[19] ),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_2/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[2] ),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_3/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[3] ),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_4/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[4] ),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_5/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[5] ),
    .X(net477));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_6/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[6] ),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_7/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[7] ),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_8/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[8] ),
    .X(net480));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y0_DSP_top/strobe_outbuf_9/_0_  (.A(\Tile_X0Y0_DSP_top/FrameStrobe_O_i[9] ),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[0] ),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[1] ),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[2] ),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[3] ),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[4] ),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[5] ),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[6] ),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[7] ),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[8] ),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/E6BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/E6BEG_i[9] ),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_0/_0_  (.A(net205),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_1/_0_  (.A(net206),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_2/_0_  (.A(net207),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_3/_0_  (.A(net208),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_4/_0_  (.A(net209),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_5/_0_  (.A(net210),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_6/_0_  (.A(net211),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_7/_0_  (.A(net212),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_8/_0_  (.A(net202),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/E6END_inbuf_9/_0_  (.A(net203),
    .X(\Tile_X0Y1_DSP_bot/E6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[0] ),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[1] ),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[10] ),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[11] ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[2] ),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[3] ),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[4] ),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[5] ),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[6] ),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[7] ),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[8] ),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/EE4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/EE4BEG_i[9] ),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_0/_0_  (.A(net223),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_1/_0_  (.A(net224),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_10/_0_  (.A(net218),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_11/_0_  (.A(net219),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_2/_0_  (.A(net225),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_3/_0_  (.A(net226),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_4/_0_  (.A(net227),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_5/_0_  (.A(net228),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_6/_0_  (.A(net214),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_7/_0_  (.A(net215),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_8/_0_  (.A(net216),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/EE4END_inbuf_9/_0_  (.A(net217),
    .X(\Tile_X0Y1_DSP_bot/EE4BEG_i[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit0  (.D(net229),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[384] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit1  (.D(net240),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[385] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit10  (.D(net230),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[394] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit11  (.D(net231),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[395] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit12  (.D(net232),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[396] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit13  (.D(net233),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[397] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit14  (.D(net234),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[398] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit15  (.D(net235),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[399] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit16  (.D(net236),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[400] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit17  (.D(net237),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[401] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit18  (.D(net238),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[402] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit19  (.D(net239),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[403] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit2  (.D(net251),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[386] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit20  (.D(net241),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[404] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit21  (.D(net242),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[405] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit22  (.D(net243),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[406] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[406] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit23  (.D(net244),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[407] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[407] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit24  (.D(net245),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[408] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[408] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit25  (.D(net246),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[409] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[409] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit26  (.D(net247),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[410] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[410] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit27  (.D(net248),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[411] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[411] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit28  (.D(net249),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[412] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[412] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit29  (.D(net250),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[413] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[413] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit3  (.D(net254),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[387] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit30  (.D(net252),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[414] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[414] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit31  (.D(net253),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[415] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[415] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit4  (.D(net255),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[388] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit5  (.D(net256),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[389] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit6  (.D(net257),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[390] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit7  (.D(net258),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[391] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit8  (.D(net259),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[392] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame0_bit9  (.D(net260),
    .GATE(net261),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[393] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit0  (.D(net229),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[64] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit1  (.D(net240),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[65] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit10  (.D(net230),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[74] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit11  (.D(net231),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[75] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit12  (.D(net232),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[76] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit13  (.D(net233),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[77] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit14  (.D(net234),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[78] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit15  (.D(net235),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[79] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit16  (.D(net236),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[80] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit17  (.D(net237),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[81] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit18  (.D(net238),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[82] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit19  (.D(net239),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[83] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit2  (.D(net251),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[66] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit20  (.D(net241),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[84] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit21  (.D(net242),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[85] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit22  (.D(net243),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[86] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit23  (.D(net244),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[87] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit24  (.D(net245),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[88] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit25  (.D(net246),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[89] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit26  (.D(net247),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[90] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit27  (.D(net248),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[91] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit28  (.D(net249),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[92] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit29  (.D(net250),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[93] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit3  (.D(net254),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[67] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit30  (.D(net252),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[94] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit31  (.D(net253),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[95] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit4  (.D(net255),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[68] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit5  (.D(net256),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[69] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit6  (.D(net257),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[70] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit7  (.D(net258),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[71] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit8  (.D(net259),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[72] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame10_bit9  (.D(net260),
    .GATE(net262),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[73] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit0  (.D(net229),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[32] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit1  (.D(net240),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[33] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit10  (.D(net230),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[42] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit11  (.D(net231),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[43] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit12  (.D(net232),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[44] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit13  (.D(net233),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[45] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit14  (.D(net234),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[46] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit15  (.D(net235),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[47] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit16  (.D(net236),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[48] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit17  (.D(net237),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[49] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit18  (.D(net238),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[50] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit19  (.D(net239),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[51] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit2  (.D(net251),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[34] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit20  (.D(net241),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[52] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit21  (.D(net242),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[53] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit22  (.D(net243),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit23  (.D(net244),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit24  (.D(net245),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[56] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit25  (.D(net246),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[57] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit26  (.D(net247),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit27  (.D(net248),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit28  (.D(net249),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[60] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit29  (.D(net250),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[61] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit3  (.D(net254),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[35] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit30  (.D(net252),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[62] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit31  (.D(net253),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[63] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit4  (.D(net255),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[36] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit5  (.D(net256),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[37] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit6  (.D(net257),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[38] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit7  (.D(net258),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[39] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit8  (.D(net259),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[40] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame11_bit9  (.D(net260),
    .GATE(net263),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[41] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit0  (.D(net229),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit1  (.D(net240),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit10  (.D(net230),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[10] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit11  (.D(net231),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[11] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit12  (.D(net232),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[12] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit13  (.D(net233),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[13] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit14  (.D(net234),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[14] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit15  (.D(net235),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[15] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit16  (.D(net236),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[16] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit17  (.D(net237),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[17] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit18  (.D(net238),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[18] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit19  (.D(net239),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[19] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit2  (.D(net251),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit20  (.D(net241),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[20] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit21  (.D(net242),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[21] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit22  (.D(net243),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[22] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit23  (.D(net244),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[23] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit24  (.D(net245),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[24] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit25  (.D(net246),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[25] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit26  (.D(net247),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[26] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit27  (.D(net248),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[27] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit28  (.D(net249),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[28] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit29  (.D(net250),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[29] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit3  (.D(net254),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit30  (.D(net252),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[30] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit31  (.D(net253),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[31] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit4  (.D(net255),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit5  (.D(net256),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit6  (.D(net257),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[6] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit7  (.D(net258),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[7] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit8  (.D(net259),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[8] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame12_bit9  (.D(net260),
    .GATE(net264),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[9] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit0  (.D(net229),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit1  (.D(net240),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit10  (.D(net230),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[362] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit11  (.D(net231),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[363] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit12  (.D(net232),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit13  (.D(net233),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit14  (.D(net234),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[366] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit15  (.D(net235),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[367] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit16  (.D(net236),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit17  (.D(net237),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit18  (.D(net238),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[370] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit19  (.D(net239),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[371] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit2  (.D(net251),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[354] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit20  (.D(net241),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit21  (.D(net242),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit22  (.D(net243),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[374] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit23  (.D(net244),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[375] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit24  (.D(net245),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit25  (.D(net246),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit26  (.D(net247),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[378] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[378] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit27  (.D(net248),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[379] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit28  (.D(net249),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit29  (.D(net250),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit3  (.D(net254),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[355] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit30  (.D(net252),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[382] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit31  (.D(net253),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[383] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit4  (.D(net255),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit5  (.D(net256),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit6  (.D(net257),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[358] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit7  (.D(net258),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[359] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit8  (.D(net259),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame1_bit9  (.D(net260),
    .GATE(net272),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit0  (.D(net229),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit1  (.D(net240),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit10  (.D(net230),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[330] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit11  (.D(net231),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[331] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit12  (.D(net232),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit13  (.D(net233),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit14  (.D(net234),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[334] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit15  (.D(net235),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[335] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit16  (.D(net236),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit17  (.D(net237),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit18  (.D(net238),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[338] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit19  (.D(net239),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[339] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit2  (.D(net251),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[322] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit20  (.D(net241),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit21  (.D(net242),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit22  (.D(net243),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[342] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit23  (.D(net244),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[343] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit24  (.D(net245),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit25  (.D(net246),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit26  (.D(net247),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[346] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit27  (.D(net248),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[347] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit28  (.D(net249),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit29  (.D(net250),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit3  (.D(net254),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[323] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit30  (.D(net252),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[350] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit31  (.D(net253),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[351] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit4  (.D(net255),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit5  (.D(net256),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit6  (.D(net257),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[326] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit7  (.D(net258),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[327] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit8  (.D(net259),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame2_bit9  (.D(net260),
    .GATE(net273),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit0  (.D(net229),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit1  (.D(net240),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit10  (.D(net230),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[298] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit11  (.D(net231),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[299] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit12  (.D(net232),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit13  (.D(net233),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit14  (.D(net234),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[302] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit15  (.D(net235),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[303] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit16  (.D(net236),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit17  (.D(net237),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit18  (.D(net238),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[306] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit19  (.D(net239),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[307] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit2  (.D(net251),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[290] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit20  (.D(net241),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit21  (.D(net242),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit22  (.D(net243),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[310] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit23  (.D(net244),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[311] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit24  (.D(net245),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit25  (.D(net246),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit26  (.D(net247),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[314] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit27  (.D(net248),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[315] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit28  (.D(net249),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit29  (.D(net250),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit3  (.D(net254),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[291] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit30  (.D(net252),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[318] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit31  (.D(net253),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[319] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit4  (.D(net255),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit5  (.D(net256),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit6  (.D(net257),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[294] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit7  (.D(net258),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[295] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit8  (.D(net259),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame3_bit9  (.D(net260),
    .GATE(net274),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit0  (.D(net229),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit1  (.D(net240),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit10  (.D(net230),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[266] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit11  (.D(net231),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[267] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit12  (.D(net232),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit13  (.D(net233),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit14  (.D(net234),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[270] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit15  (.D(net235),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[271] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit16  (.D(net236),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit17  (.D(net237),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit18  (.D(net238),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[274] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit19  (.D(net239),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[275] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit2  (.D(net251),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[258] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit20  (.D(net241),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit21  (.D(net242),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit22  (.D(net243),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[278] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit23  (.D(net244),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[279] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit24  (.D(net245),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit25  (.D(net246),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit26  (.D(net247),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[282] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit27  (.D(net248),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[283] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit28  (.D(net249),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit29  (.D(net250),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit3  (.D(net254),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[259] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit30  (.D(net252),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[286] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit31  (.D(net253),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[287] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit4  (.D(net255),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit5  (.D(net256),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit6  (.D(net257),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[262] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit7  (.D(net258),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[263] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit8  (.D(net259),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame4_bit9  (.D(net260),
    .GATE(net275),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit0  (.D(net229),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[224] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit1  (.D(net240),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[225] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit10  (.D(net230),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[234] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit11  (.D(net231),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[235] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit12  (.D(net232),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[236] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit13  (.D(net233),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[237] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit14  (.D(net234),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[238] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit15  (.D(net235),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[239] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit16  (.D(net236),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[240] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit17  (.D(net237),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[241] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit18  (.D(net238),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[242] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit19  (.D(net239),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[243] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit2  (.D(net251),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[226] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit20  (.D(net241),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[244] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit21  (.D(net242),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[245] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit22  (.D(net243),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[246] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit23  (.D(net244),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[247] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit24  (.D(net245),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[248] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit25  (.D(net246),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[249] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit26  (.D(net247),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[250] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit27  (.D(net248),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[251] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit28  (.D(net249),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[252] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit29  (.D(net250),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[253] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit3  (.D(net254),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[227] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit30  (.D(net252),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[254] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit31  (.D(net253),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[255] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit4  (.D(net255),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[228] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit5  (.D(net256),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[229] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit6  (.D(net257),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[230] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit7  (.D(net258),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[231] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit8  (.D(net259),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[232] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame5_bit9  (.D(net260),
    .GATE(net276),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[233] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit0  (.D(net229),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[192] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit1  (.D(net240),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[193] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit10  (.D(net230),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[202] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit11  (.D(net231),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[203] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit12  (.D(net232),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[204] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit13  (.D(net233),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[205] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit14  (.D(net234),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[206] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit15  (.D(net235),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[207] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit16  (.D(net236),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[208] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit17  (.D(net237),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[209] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit18  (.D(net238),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[210] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit19  (.D(net239),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[211] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit2  (.D(net251),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[194] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit20  (.D(net241),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[212] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit21  (.D(net242),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[213] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit22  (.D(net243),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[214] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit23  (.D(net244),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[215] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit24  (.D(net245),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[216] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit25  (.D(net246),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[217] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit26  (.D(net247),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[218] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit27  (.D(net248),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[219] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit28  (.D(net249),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[220] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit29  (.D(net250),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[221] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit3  (.D(net254),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[195] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit30  (.D(net252),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[222] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit31  (.D(net253),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[223] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit4  (.D(net255),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[196] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit5  (.D(net256),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[197] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit6  (.D(net257),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[198] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit7  (.D(net258),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[199] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit8  (.D(net259),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[200] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame6_bit9  (.D(net260),
    .GATE(net277),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[201] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit0  (.D(net229),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[160] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit1  (.D(net240),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[161] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit10  (.D(net230),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[170] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit11  (.D(net231),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[171] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit12  (.D(net232),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[172] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit13  (.D(net233),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[173] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit14  (.D(net234),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[174] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit15  (.D(net235),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[175] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit16  (.D(net236),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[176] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit17  (.D(net237),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[177] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit18  (.D(net238),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[178] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit19  (.D(net239),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[179] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit2  (.D(net251),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[162] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit20  (.D(net241),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[180] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit21  (.D(net242),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[181] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit22  (.D(net243),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[182] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit23  (.D(net244),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[183] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit24  (.D(net245),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[184] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit25  (.D(net246),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[185] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit26  (.D(net247),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[186] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit27  (.D(net248),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[187] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit28  (.D(net249),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[188] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit29  (.D(net250),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[189] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit3  (.D(net254),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[163] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit30  (.D(net252),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[190] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit31  (.D(net253),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[191] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit4  (.D(net255),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[164] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit5  (.D(net256),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[165] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit6  (.D(net257),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[166] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit7  (.D(net258),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[167] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit8  (.D(net259),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[168] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame7_bit9  (.D(net260),
    .GATE(net278),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[169] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit0  (.D(net229),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[128] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit1  (.D(net240),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[129] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit10  (.D(net230),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[138] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit11  (.D(net231),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[139] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit12  (.D(net232),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[140] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit13  (.D(net233),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[141] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit14  (.D(net234),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[142] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit15  (.D(net235),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[143] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit16  (.D(net236),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[144] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit17  (.D(net237),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[145] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit18  (.D(net238),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[146] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit19  (.D(net239),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[147] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit2  (.D(net251),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[130] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit20  (.D(net241),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[148] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit21  (.D(net242),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[149] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit22  (.D(net243),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[150] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit23  (.D(net244),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[151] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit24  (.D(net245),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[152] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit25  (.D(net246),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[153] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit26  (.D(net247),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[154] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit27  (.D(net248),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[155] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit28  (.D(net249),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit29  (.D(net250),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit3  (.D(net254),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[131] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit30  (.D(net252),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[158] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit31  (.D(net253),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[159] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit4  (.D(net255),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[132] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit5  (.D(net256),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[133] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit6  (.D(net257),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[134] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit7  (.D(net258),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[135] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit8  (.D(net259),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[136] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame8_bit9  (.D(net260),
    .GATE(net279),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[137] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit0  (.D(net229),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[96] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit1  (.D(net240),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[97] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit10  (.D(net230),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[106] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit11  (.D(net231),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[107] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit12  (.D(net232),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[108] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit13  (.D(net233),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[109] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit14  (.D(net234),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit15  (.D(net235),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit16  (.D(net236),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[112] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit17  (.D(net237),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[113] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit18  (.D(net238),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit19  (.D(net239),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit2  (.D(net251),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[98] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit20  (.D(net241),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[116] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit21  (.D(net242),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[117] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit22  (.D(net243),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[118] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit23  (.D(net244),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[119] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit24  (.D(net245),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[120] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit25  (.D(net246),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[121] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit26  (.D(net247),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[122] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit27  (.D(net248),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[123] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit28  (.D(net249),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[124] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit29  (.D(net250),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[125] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit3  (.D(net254),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[99] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit30  (.D(net252),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[126] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit31  (.D(net253),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[127] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit4  (.D(net255),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[100] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit5  (.D(net256),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[101] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit6  (.D(net257),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[102] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit7  (.D(net258),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[103] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit8  (.D(net259),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[104] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_ConfigMem/Inst_frame9_bit9  (.D(net260),
    .GATE(net280),
    .Q(\Tile_X0Y1_DSP_bot/ConfigBits[105] ),
    .Q_N(\Tile_X0Y1_DSP_bot/ConfigBits_N[105] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_04_  (.A(\Tile_X0Y0_top2bot[0] ),
    .X(\Tile_X0Y1_DSP_bot/A4 ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_05_  (.A(\Tile_X0Y0_top2bot[1] ),
    .X(\Tile_X0Y1_DSP_bot/A5 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_06_  (.A(\Tile_X0Y0_top2bot[2] ),
    .X(\Tile_X0Y1_DSP_bot/A6 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_07_  (.A(\Tile_X0Y0_top2bot[3] ),
    .X(\Tile_X0Y1_DSP_bot/A7 ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_08_  (.A(\Tile_X0Y0_top2bot[4] ),
    .X(\Tile_X0Y1_DSP_bot/B4 ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_09_  (.A(\Tile_X0Y0_top2bot[5] ),
    .X(\Tile_X0Y1_DSP_bot/B5 ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_10_  (.A(\Tile_X0Y0_top2bot[6] ),
    .X(\Tile_X0Y1_DSP_bot/B6 ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_11_  (.A(\Tile_X0Y0_top2bot[7] ),
    .X(\Tile_X0Y1_DSP_bot/B7 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_12_  (.A(\Tile_X0Y0_top2bot[8] ),
    .X(\Tile_X0Y1_DSP_bot/C10 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_13_  (.A(\Tile_X0Y0_top2bot[9] ),
    .X(\Tile_X0Y1_DSP_bot/C11 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_14_  (.A(\Tile_X0Y0_top2bot[10] ),
    .X(\Tile_X0Y1_DSP_bot/C12 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_15_  (.A(\Tile_X0Y0_top2bot[11] ),
    .X(\Tile_X0Y1_DSP_bot/C13 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_16_  (.A(\Tile_X0Y0_top2bot[12] ),
    .X(\Tile_X0Y1_DSP_bot/C14 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_17_  (.A(\Tile_X0Y0_top2bot[13] ),
    .X(\Tile_X0Y1_DSP_bot/C15 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_18_  (.A(\Tile_X0Y0_top2bot[14] ),
    .X(\Tile_X0Y1_DSP_bot/C16 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_19_  (.A(\Tile_X0Y0_top2bot[15] ),
    .X(\Tile_X0Y1_DSP_bot/C17 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_20_  (.A(\Tile_X0Y0_top2bot[16] ),
    .X(\Tile_X0Y1_DSP_bot/C18 ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_21_  (.A(\Tile_X0Y0_top2bot[17] ),
    .X(\Tile_X0Y1_DSP_bot/C19 ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_22_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[0] ),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_23_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[1] ),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_24_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_25_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_26_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_27_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[5] ),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_28_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_29_  (.A(\Tile_X0Y1_DSP_bot/JE2BEG[7] ),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_30_  (.A(net193),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_31_  (.A(net194),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_32_  (.A(net195),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_33_  (.A(net196),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_34_  (.A(net197),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_35_  (.A(net198),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_36_  (.A(net199),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_37_  (.A(net200),
    .X(net602));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_38_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[0] ),
    .X(\Tile_X0Y1_N2BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_39_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[1] ),
    .X(\Tile_X0Y1_N2BEG[1] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_40_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .X(\Tile_X0Y1_N2BEG[2] ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_41_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .X(\Tile_X0Y1_N2BEG[3] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_42_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .X(\Tile_X0Y1_N2BEG[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_43_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[5] ),
    .X(\Tile_X0Y1_N2BEG[5] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_44_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[6] ),
    .X(\Tile_X0Y1_N2BEG[6] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_45_  (.A(\Tile_X0Y1_DSP_bot/JN2BEG[7] ),
    .X(\Tile_X0Y1_N2BEG[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_46_  (.A(net293),
    .X(\Tile_X0Y1_N2BEGb[0] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_47_  (.A(net294),
    .X(\Tile_X0Y1_N2BEGb[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_48_  (.A(net295),
    .X(\Tile_X0Y1_N2BEGb[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_49_  (.A(net296),
    .X(\Tile_X0Y1_N2BEGb[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_50_  (.A(net297),
    .X(\Tile_X0Y1_N2BEGb[4] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_51_  (.A(net298),
    .X(\Tile_X0Y1_N2BEGb[5] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_52_  (.A(net299),
    .X(\Tile_X0Y1_N2BEGb[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_53_  (.A(net300),
    .X(\Tile_X0Y1_N2BEGb[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_54_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[0] ),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_55_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[1] ),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_56_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_57_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_58_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_59_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[5] ),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_60_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[6] ),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_61_  (.A(\Tile_X0Y1_DSP_bot/JS2BEG[7] ),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_62_  (.A(\Tile_X0Y0_S2BEG[0] ),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_63_  (.A(\Tile_X0Y0_S2BEG[1] ),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_64_  (.A(\Tile_X0Y0_S2BEG[2] ),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_65_  (.A(\Tile_X0Y0_S2BEG[3] ),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_66_  (.A(\Tile_X0Y0_S2BEG[4] ),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_67_  (.A(\Tile_X0Y0_S2BEG[5] ),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_68_  (.A(\Tile_X0Y0_S2BEG[6] ),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_69_  (.A(\Tile_X0Y0_S2BEG[7] ),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_70_  (.A(net338),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_71_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[1] ),
    .X(net720));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_72_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_73_  (.A(net341),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_74_  (.A(net342),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_75_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_76_  (.A(\Tile_X0Y1_DSP_bot/JW2BEG[6] ),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_77_  (.A(net345),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_78_  (.A(net346),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_79_  (.A(net347),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_80_  (.A(net348),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_81_  (.A(net349),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_82_  (.A(net350),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_83_  (.A(net351),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_84_  (.A(net352),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_85_  (.A(net353),
    .X(net734));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_86_  (.A(\Tile_X0Y1_DSP_bot/Q10 ),
    .X(\Tile_X0Y1_bot2top[0] ));
 sky130_fd_sc_hd__clkbuf_16 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_87_  (.A(\Tile_X0Y1_DSP_bot/Q11 ),
    .X(\Tile_X0Y1_bot2top[1] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_88_  (.A(\Tile_X0Y1_DSP_bot/Q12 ),
    .X(\Tile_X0Y1_bot2top[2] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_89_  (.A(\Tile_X0Y1_DSP_bot/Q13 ),
    .X(\Tile_X0Y1_bot2top[3] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_90_  (.A(\Tile_X0Y1_DSP_bot/Q14 ),
    .X(\Tile_X0Y1_bot2top[4] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_91_  (.A(\Tile_X0Y1_DSP_bot/Q15 ),
    .X(\Tile_X0Y1_bot2top[5] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_92_  (.A(\Tile_X0Y1_DSP_bot/Q16 ),
    .X(\Tile_X0Y1_bot2top[6] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_93_  (.A(\Tile_X0Y1_DSP_bot/Q17 ),
    .X(\Tile_X0Y1_bot2top[7] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_94_  (.A(\Tile_X0Y1_DSP_bot/Q18 ),
    .X(\Tile_X0Y1_bot2top[8] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/_95_  (.A(\Tile_X0Y1_DSP_bot/Q19 ),
    .X(\Tile_X0Y1_bot2top[9] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0  (.A0(net184),
    .A1(net337),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(\Tile_X0Y1_DSP_bot/Q1 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[54] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[55] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[56] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[57] ),
    .X(net604));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0  (.A0(net183),
    .A1(net336),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(\Tile_X0Y1_DSP_bot/Q1 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[58] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[59] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[60] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[61] ),
    .X(net605));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net286),
    .A2(net308),
    .A3(net220),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q1 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[288] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[289] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[290] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[291] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net287),
    .A2(net309),
    .A3(net187),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[2] ),
    .A2(net340),
    .A3(net375),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[292] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[293] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[294] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[295] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net288),
    .A2(net310),
    .A3(net188),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[3] ),
    .A2(net341),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[296] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[297] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[298] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[299] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net289),
    .A2(net301),
    .A3(net189),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[4] ),
    .A2(net342),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[300] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[301] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[302] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[303] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[5] ),
    .A3(net335),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[304] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[305] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[306] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[307] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_S2BEGb[6] ),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[308] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[309] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[310] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[311] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[312] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[313] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[314] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[315] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net185),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_SS4BEG[0] ),
    .A3(net366),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[316] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[317] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[318] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[319] ),
    .X(\Tile_X0Y1_DSP_bot/JE2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0  (.A0(net286),
    .A1(net308),
    .A2(net184),
    .A3(net186),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_SS4BEG[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2  (.A0(net764),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[256] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[257] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[258] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[259] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0  (.A0(net287),
    .A1(net309),
    .A2(net181),
    .A3(net187),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[2] ),
    .A2(net340),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[260] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[261] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[262] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[263] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0  (.A0(net288),
    .A1(net310),
    .A2(net182),
    .A3(net188),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[3] ),
    .A2(net341),
    .A3(net373),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[264] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[265] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[266] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[267] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0  (.A0(net289),
    .A1(net301),
    .A2(net183),
    .A3(net189),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[4] ),
    .A2(net342),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[268] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[269] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[270] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[271] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S2BEGb[5] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[272] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[273] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[274] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[275] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[2] ),
    .A1(\Tile_X0Y0_S2BEGb[6] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[276] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[277] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[278] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[279] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[3] ),
    .A1(\Tile_X0Y0_S2BEGb[7] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[280] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[281] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[282] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[283] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net213),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S2BEGb[0] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[284] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[285] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[286] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[287] ),
    .X(\Tile_X0Y1_DSP_bot/JN2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0  (.A0(net324),
    .A1(net184),
    .A2(net186),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[1] ),
    .A1(\Tile_X0Y0_S4BEG[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q1 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[320] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[321] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[322] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[323] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0  (.A0(net325),
    .A1(net181),
    .A2(net221),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S4BEG[2] ),
    .A1(\Tile_X0Y0_SS4BEG[2] ),
    .A2(net340),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[324] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[325] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[326] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[327] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0  (.A0(net326),
    .A1(net182),
    .A2(net188),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[3] ),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net341),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[328] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[329] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[330] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[331] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0  (.A0(net289),
    .A1(net183),
    .A2(net189),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[4] ),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net342),
    .A3(net374),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[332] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[333] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[334] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[335] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S2BEGb[5] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[336] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[337] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[338] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[339] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[2] ),
    .A1(\Tile_X0Y0_S2BEGb[6] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[340] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[341] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[342] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[343] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[3] ),
    .A1(\Tile_X0Y0_S2BEGb[7] ),
    .A2(net335),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[344] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[345] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[346] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[347] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net185),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S2BEGb[0] ),
    .A2(net334),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[348] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[349] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[350] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[351] ),
    .X(\Tile_X0Y1_DSP_bot/JS2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net286),
    .A2(net186),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[1] ),
    .A1(\Tile_X0Y0_S4BEG[1] ),
    .A2(net339),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q1 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[352] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[353] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[354] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[355] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net287),
    .A2(net187),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[2] ),
    .A1(\Tile_X0Y0_S4BEG[2] ),
    .A2(net340),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q2 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[356] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[357] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[358] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[359] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net288),
    .A2(net188),
    .A3(net204),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[3] ),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net341),
    .A3(net357),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q3 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(net763),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[360] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[361] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[362] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[363] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net289),
    .A2(net189),
    .A3(net201),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S2BEGb[4] ),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net342),
    .A3(net354),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[364] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[365] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[366] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[367] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net290),
    .A2(net182),
    .A3(net190),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[5] ),
    .A3(net335),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[368] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[369] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[370] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[371] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net291),
    .A2(net183),
    .A3(net191),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_S2BEGb[6] ),
    .A3(net336),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q6 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[372] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[373] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[374] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[375] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net292),
    .A2(net184),
    .A3(net192),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[1] ),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net337),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(net764),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(\Tile_X0Y1_DSP_bot/Q7 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[376] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[377] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[378] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[379] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net285),
    .A2(net181),
    .A3(net185),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1  (.A0(\Tile_X0Y0_S1BEG[0] ),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(\Tile_X0Y0_S2BEGb[0] ),
    .A3(net334),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/Q1 ),
    .A2(\Tile_X0Y1_DSP_bot/Q2 ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/Q5 ),
    .A2(net763),
    .A3(\Tile_X0Y1_DSP_bot/Q8 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[380] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[381] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[382] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[383] ),
    .X(\Tile_X0Y1_DSP_bot/JW2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0  (.A0(net184),
    .A1(net337),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(net764),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q6 ),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[110] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[111] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[112] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[113] ),
    .X(net736));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0  (.A0(net183),
    .A1(net336),
    .A2(\Tile_X0Y1_DSP_bot/Q0 ),
    .A3(net764),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/Q3 ),
    .A2(\Tile_X0Y1_DSP_bot/Q4 ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/Q6 ),
    .A1(\Tile_X0Y1_DSP_bot/Q7 ),
    .A2(\Tile_X0Y1_DSP_bot/Q8 ),
    .A3(\Tile_X0Y1_DSP_bot/Q9 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[114] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[115] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[116] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[117] ),
    .X(net737));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst0  (.A0(net299),
    .A1(net193),
    .A2(net199),
    .A3(\Tile_X0Y0_S2BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst1  (.A0(net346),
    .A1(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst2  (.A0(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst3  (.A0(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .A2(net765),
    .A3(net766),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[156] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[157] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__conb_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst3_765  (.LO(net765));
 sky130_fd_sc_hd__conb_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst3_766  (.HI(net766));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_inst4  (.A0(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out1 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out2 ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux161_buf_clr/cus_mux41_buf_out3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[158] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[159] ),
    .X(\Tile_X0Y1_DSP_bot/clr ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A0  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[118] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[119] ),
    .X(\Tile_X0Y1_DSP_bot/A0 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A1  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[120] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[121] ),
    .X(\Tile_X0Y1_DSP_bot/A1 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A2  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[122] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[123] ),
    .X(\Tile_X0Y1_DSP_bot/A2 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_A3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[124] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[125] ),
    .X(\Tile_X0Y1_DSP_bot/A3 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B0  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[126] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[127] ),
    .X(\Tile_X0Y1_DSP_bot/B0 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B1  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[128] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[129] ),
    .X(\Tile_X0Y1_DSP_bot/B1 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B2  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[130] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[131] ),
    .X(\Tile_X0Y1_DSP_bot/B2 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_B3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[132] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[133] ),
    .X(\Tile_X0Y1_DSP_bot/B3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C0  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[134] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[135] ),
    .X(\Tile_X0Y1_DSP_bot/C0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C1  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[136] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[137] ),
    .X(\Tile_X0Y1_DSP_bot/C1 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C2  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[138] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[139] ),
    .X(\Tile_X0Y1_DSP_bot/C2 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C3  (.A0(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[140] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[141] ),
    .X(\Tile_X0Y1_DSP_bot/C3 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C4  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[0] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[142] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[143] ),
    .X(\Tile_X0Y1_DSP_bot/C4 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C5  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[1] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[144] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[145] ),
    .X(\Tile_X0Y1_DSP_bot/C5 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C6  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[146] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[147] ),
    .X(\Tile_X0Y1_DSP_bot/C6 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_C7  (.A0(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[3] ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[148] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[149] ),
    .X(\Tile_X0Y1_DSP_bot/C7 ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q3 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[34] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[35] ),
    .X(net583));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG1  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[36] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[37] ),
    .X(net584));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG2  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[38] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[39] ),
    .X(net585));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_E1BEG3  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[40] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[41] ),
    .X(net586));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(net291),
    .A1(net191),
    .A2(\Tile_X0Y0_SS4BEG[3] ),
    .A3(net344),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[224] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[225] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(net317),
    .A1(net187),
    .A2(\Tile_X0Y0_S2BEGb[2] ),
    .A3(net340),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[226] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[227] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(net289),
    .A1(net213),
    .A2(\Tile_X0Y0_S2BEGb[4] ),
    .A3(net342),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[228] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[229] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(net285),
    .A1(net185),
    .A2(\Tile_X0Y0_S2BEGb[0] ),
    .A3(net375),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[230] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[231] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(net326),
    .A1(net191),
    .A2(\Tile_X0Y0_S2BEGb[6] ),
    .A3(net344),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[232] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[233] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(net287),
    .A1(net187),
    .A2(\Tile_X0Y0_S2BEGb[2] ),
    .A3(net374),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[234] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[235] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(net289),
    .A1(net189),
    .A2(\Tile_X0Y0_SS4BEG[2] ),
    .A3(net342),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[236] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[237] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(net285),
    .A1(net220),
    .A2(\Tile_X0Y0_S2BEGb[0] ),
    .A3(net338),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[238] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[239] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(net292),
    .A1(net221),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net345),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[240] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[241] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(net288),
    .A1(net188),
    .A2(\Tile_X0Y0_S2BEGb[3] ),
    .A3(net373),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[242] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[243] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(net290),
    .A1(net190),
    .A2(\Tile_X0Y0_SS4BEG[1] ),
    .A3(net343),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[244] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[245] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(net325),
    .A1(net186),
    .A2(\Tile_X0Y0_S2BEGb[1] ),
    .A3(net339),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[246] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[247] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(net292),
    .A1(net192),
    .A2(\Tile_X0Y0_S2BEGb[7] ),
    .A3(net366),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[248] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[249] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(net288),
    .A1(net188),
    .A2(\Tile_X0Y0_SS4BEG[0] ),
    .A3(net341),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[250] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[251] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(net324),
    .A1(net190),
    .A2(\Tile_X0Y0_S2BEGb[5] ),
    .A3(net343),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[252] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[253] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(net286),
    .A1(net222),
    .A2(\Tile_X0Y0_S2BEGb[1] ),
    .A3(net339),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[254] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[255] ),
    .X(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(net299),
    .A1(\Tile_X0Y0_S2BEG[6] ),
    .A2(net352),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[160] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[161] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net195),
    .A1(\Tile_X0Y0_S2BEG[2] ),
    .A2(net348),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[162] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[163] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(net297),
    .A1(net197),
    .A2(net350),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[164] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[165] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(net293),
    .A1(net193),
    .A2(\Tile_X0Y0_S2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[166] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[167] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[192] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[193] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[194] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[195] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[196] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[197] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[198] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[199] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net199),
    .A1(\Tile_X0Y0_S2BEG[6] ),
    .A2(net352),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[168] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[169] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(net295),
    .A1(net195),
    .A2(net348),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[170] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[171] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(net297),
    .A1(net197),
    .A2(\Tile_X0Y0_S2BEG[4] ),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[172] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[173] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(net293),
    .A1(\Tile_X0Y0_S2BEG[0] ),
    .A2(net346),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[174] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[175] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[200] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[201] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[202] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[203] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[204] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[205] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[206] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[207] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(net299),
    .A1(net199),
    .A2(net352),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[176] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[177] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(net295),
    .A1(net195),
    .A2(\Tile_X0Y0_S2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[178] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[179] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(net297),
    .A1(\Tile_X0Y0_S2BEG[4] ),
    .A2(net350),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[180] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[181] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net193),
    .A1(\Tile_X0Y0_S2BEG[0] ),
    .A2(net346),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[182] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[183] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[208] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[209] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[210] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[211] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[212] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[213] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[214] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[215] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(net299),
    .A1(net199),
    .A2(\Tile_X0Y0_S2BEG[6] ),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[184] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[185] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(net295),
    .A1(\Tile_X0Y0_S2BEG[2] ),
    .A2(net348),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[186] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[187] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net197),
    .A1(\Tile_X0Y0_S2BEG[4] ),
    .A2(net350),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[188] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[189] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(net293),
    .A1(net193),
    .A2(net346),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[190] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[191] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(net300),
    .A1(net200),
    .A2(\Tile_X0Y0_S2BEG[7] ),
    .A3(net353),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[216] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[217] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(net296),
    .A1(net196),
    .A2(\Tile_X0Y0_S2BEG[3] ),
    .A3(net349),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[218] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[219] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(net298),
    .A1(net198),
    .A2(\Tile_X0Y0_S2BEG[5] ),
    .A3(net351),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[220] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[221] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(net294),
    .A1(net194),
    .A2(\Tile_X0Y0_S2BEG[1] ),
    .A3(net347),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[222] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[223] ),
    .X(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(net326),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net366),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[384] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[385] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net221),
    .A1(\Tile_X0Y0_S4BEG[2] ),
    .A2(net345),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[386] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[387] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(net308),
    .A1(net204),
    .A2(net357),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[388] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[389] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(net301),
    .A1(net201),
    .A2(\Tile_X0Y0_S4BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[390] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[391] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net188),
    .A1(\Tile_X0Y0_SS4BEG[3] ),
    .A2(net374),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[392] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[393] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(net309),
    .A1(net187),
    .A2(net345),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[394] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[395] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(net324),
    .A1(net220),
    .A2(\Tile_X0Y0_S4BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[396] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[397] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(net301),
    .A1(\Tile_X0Y0_SS4BEG[0] ),
    .A2(net354),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[398] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[399] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(net310),
    .A1(net188),
    .A2(net341),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[400] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[401] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(net325),
    .A1(net187),
    .A2(\Tile_X0Y0_S4BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[402] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[403] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(net308),
    .A1(\Tile_X0Y0_SS4BEG[1] ),
    .A2(net342),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[404] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[405] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net222),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net373),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[406] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[407] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(net310),
    .A1(net213),
    .A2(\Tile_X0Y0_S4BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[408] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[409] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(net309),
    .A1(\Tile_X0Y0_SS4BEG[2] ),
    .A2(net340),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[410] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[411] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net204),
    .A1(\Tile_X0Y0_S4BEG[1] ),
    .A2(net375),
    .A3(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[412] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[413] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(net317),
    .A1(net201),
    .A2(net338),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[4] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[414] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[415] ),
    .X(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q2 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[6] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[7] ),
    .X(\Tile_X0Y1_N1BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(\Tile_X0Y1_DSP_bot/Q3 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[8] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[9] ),
    .X(\Tile_X0Y1_N1BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[10] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[11] ),
    .X(\Tile_X0Y1_N1BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[12] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[13] ),
    .X(\Tile_X0Y1_N1BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG0  (.A0(net287),
    .A1(net308),
    .A2(net204),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[14] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[15] ),
    .X(\Tile_X0Y1_N4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG1  (.A0(net288),
    .A1(net309),
    .A2(net201),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[16] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[17] ),
    .X(\Tile_X0Y1_N4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG2  (.A0(net285),
    .A1(net310),
    .A2(net357),
    .A3(\Tile_X0Y1_DSP_bot/Q6 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[18] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[19] ),
    .X(\Tile_X0Y1_N4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_N4BEG3  (.A0(net286),
    .A1(net301),
    .A2(net354),
    .A3(\Tile_X0Y1_DSP_bot/Q7 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[20] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[21] ),
    .X(\Tile_X0Y1_N4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q4 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[62] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[63] ),
    .X(net663));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[64] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[65] ),
    .X(net664));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[66] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[67] ),
    .X(net665));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[68] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[69] ),
    .X(net666));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG0  (.A0(net204),
    .A1(\Tile_X0Y0_S2BEGb[2] ),
    .A2(\Tile_X0Y0_S4BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/Q0 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[70] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[71] ),
    .X(net686));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG1  (.A0(net201),
    .A1(\Tile_X0Y0_S2BEGb[3] ),
    .A2(\Tile_X0Y0_S4BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/Q1 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[72] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[73] ),
    .X(net687));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG2  (.A0(\Tile_X0Y0_S2BEGb[0] ),
    .A1(\Tile_X0Y0_S4BEG[3] ),
    .A2(net357),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[74] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[75] ),
    .X(net688));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_S4BEG3  (.A0(\Tile_X0Y0_S2BEGb[1] ),
    .A1(\Tile_X0Y0_S4BEG[0] ),
    .A2(net354),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[76] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[77] ),
    .X(net689));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(\Tile_X0Y1_DSP_bot/Q5 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[3] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[90] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[91] ),
    .X(net715));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[0] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[92] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[93] ),
    .X(net716));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[94] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[95] ),
    .X(net717));
 sky130_fd_sc_hd__mux4_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(\Tile_X0Y1_DSP_bot/Q0 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/JS2BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J_l_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[96] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[97] ),
    .X(net718));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_DSP_bot/JN2BEG[4] ),
    .A1(\Tile_X0Y1_DSP_bot/JN2BEG[6] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[4] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[150] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[151] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/JS2BEG[4] ),
    .A1(\Tile_X0Y1_DSP_bot/JS2BEG[6] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[4] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[6] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[150] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[151] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[152] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[152] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C8/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y1_DSP_bot/C8 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_inst0  (.A0(\Tile_X0Y1_DSP_bot/JN2BEG[5] ),
    .A1(\Tile_X0Y1_DSP_bot/JN2BEG[7] ),
    .A2(\Tile_X0Y1_DSP_bot/JE2BEG[5] ),
    .A3(\Tile_X0Y1_DSP_bot/JE2BEG[7] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[153] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[154] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/JS2BEG[5] ),
    .A1(\Tile_X0Y1_DSP_bot/JS2BEG[7] ),
    .A2(\Tile_X0Y1_DSP_bot/JW2BEG[5] ),
    .A3(\Tile_X0Y1_DSP_bot/JW2BEG[7] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[153] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[154] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[155] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[155] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_C9/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y1_DSP_bot/C9 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net183),
    .A2(\Tile_X0Y0_S1BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[42] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[43] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[42] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[43] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[44] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[44] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_1_ ),
    .Y(net618));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net184),
    .A2(\Tile_X0Y0_S1BEG[3] ),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[45] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[46] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[45] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[46] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[47] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[47] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_1_ ),
    .Y(net619));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net181),
    .A2(\Tile_X0Y0_S1BEG[0] ),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[48] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[49] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[48] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[49] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[50] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[50] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_1_ ),
    .Y(net620));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net182),
    .A2(\Tile_X0Y0_S1BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[51] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[52] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[0] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[51] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[52] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[53] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[53] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_1_ ),
    .Y(net621));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net183),
    .A2(net336),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[22] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[23] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[22] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[23] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[24] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[24] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y1_NN4BEG[12] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net184),
    .A2(net337),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[25] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[26] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[25] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[26] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[27] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[27] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y1_NN4BEG[13] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net181),
    .A2(net334),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[28] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[29] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[28] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[29] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[30] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[30] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y1_NN4BEG[14] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net182),
    .A2(net335),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[31] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[32] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[1] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[31] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[32] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[33] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[33] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_1_ ),
    .Y(\Tile_X0Y1_NN4BEG[15] ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(net183),
    .A2(net336),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[78] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[79] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1  (.A0(net763),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[78] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[79] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[80] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[80] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_1_ ),
    .Y(net702));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(net184),
    .A2(net337),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[81] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[82] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[81] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[82] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[83] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[83] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_1_ ),
    .Y(net703));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(net181),
    .A2(net334),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[84] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[85] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[84] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[85] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[86] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[86] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_1_ ),
    .Y(net704));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(net182),
    .A2(net335),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[87] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[88] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[3] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[87] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[88] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[89] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[89] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_1_ ),
    .Y(net705));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0  (.A0(net283),
    .A1(\Tile_X0Y0_S1BEG[2] ),
    .A2(net336),
    .A3(\Tile_X0Y1_DSP_bot/Q2 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[98] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[99] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q6 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_GH_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[98] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[99] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[100] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[100] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_1_ ),
    .Y(net750));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0  (.A0(net284),
    .A1(\Tile_X0Y0_S1BEG[3] ),
    .A2(net337),
    .A3(\Tile_X0Y1_DSP_bot/Q3 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[101] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[102] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q7 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_ABa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_CDa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_EF_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[101] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[102] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[103] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[103] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_1_ ),
    .Y(net751));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0  (.A0(net281),
    .A1(\Tile_X0Y0_S1BEG[0] ),
    .A2(net334),
    .A3(\Tile_X0Y1_DSP_bot/Q4 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[104] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[105] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q8 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFb_BEG[1] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHb_BEG[1] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_CD_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[104] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[105] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[106] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[106] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_1_ ),
    .Y(net752));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0  (.A0(net282),
    .A1(\Tile_X0Y0_S1BEG[1] ),
    .A2(net335),
    .A3(\Tile_X0Y1_DSP_bot/Q5 ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[107] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[108] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1  (.A0(\Tile_X0Y1_DSP_bot/Q9 ),
    .A1(\Tile_X0Y1_DSP_bot/J2MID_EFa_BEG[2] ),
    .A2(\Tile_X0Y1_DSP_bot/J2MID_GHa_BEG[2] ),
    .A3(\Tile_X0Y1_DSP_bot/J2END_AB_BEG[2] ),
    .S0(\Tile_X0Y1_DSP_bot/ConfigBits[107] ),
    .S1(\Tile_X0Y1_DSP_bot/ConfigBits[108] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_2_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_3_  (.A(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[109] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_4_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[109] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_DSP_bot_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_1_ ),
    .Y(net753));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0843_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0844_  (.A0(\Tile_X0Y1_DSP_bot/C0 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[0] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0022_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0845_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0022_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0846_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0847_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0848_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0849_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[0] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0850_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0851_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0852_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[0] ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0853_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .B_N(\Tile_X0Y1_DSP_bot/B0 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ));
 sky130_fd_sc_hd__nand2_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0854_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0855_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0856_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0857_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0023_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0858_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0036_ ));
 sky130_fd_sc_hd__a21bo_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0859_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0036_ ),
    .X(\Tile_X0Y1_DSP_bot/Q0 ));
 sky130_fd_sc_hd__buf_6 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0860_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0861_  (.A(\Tile_X0Y1_DSP_bot/A1 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0862_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0863_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0864_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0865_  (.A(\Tile_X0Y1_DSP_bot/B1 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0042_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0866_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[1] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0867_  (.A1(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0042_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0868_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0869_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0870_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0871_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .A2(\Tile_X0Y1_DSP_bot/B0 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0872_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0039_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0873_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .A2(\Tile_X0Y1_DSP_bot/B1 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0043_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0874_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ));
 sky130_fd_sc_hd__or4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0875_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0876_  (.A0(\Tile_X0Y1_DSP_bot/C1 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[1] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0053_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0877_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0053_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0878_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0055_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0879_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0056_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0880_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0055_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0056_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ));
 sky130_fd_sc_hd__xnor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0881_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0882_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0059_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0883_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0059_ ),
    .Y(\Tile_X0Y1_DSP_bot/Q1 ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0884_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0046_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0054_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0057_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0885_  (.A(\Tile_X0Y1_DSP_bot/A2 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0886_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[2] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0887_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ));
 sky130_fd_sc_hd__and2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0888_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ));
 sky130_fd_sc_hd__nor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0889_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0038_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0890_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0891_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0892_  (.A(\Tile_X0Y1_DSP_bot/B2 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0893_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0894_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0895_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0896_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0897_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0061_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0062_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0898_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0899_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0900_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ));
 sky130_fd_sc_hd__o311a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0901_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0902_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0078_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0903_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[1] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ));
 sky130_fd_sc_hd__o21a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0904_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0068_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0069_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ));
 sky130_fd_sc_hd__o2bb2a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0905_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0078_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ));
 sky130_fd_sc_hd__nor3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0906_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0907_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0077_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0081_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0052_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0083_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0908_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0083_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0909_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[3] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0910_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[2] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0911_  (.A0(\Tile_X0Y1_DSP_bot/C2 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[2] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0087_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0912_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0088_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0913_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0087_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0088_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0914_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0915_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0084_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0089_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0916_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0092_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0917_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0092_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0918_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0919_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0095_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0920_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0095_ ),
    .X(\Tile_X0Y1_DSP_bot/Q2 ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0921_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[3] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0096_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0922_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .A2(\Tile_X0Y1_DSP_bot/C3 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0096_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0923_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0924_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0925_  (.A(\Tile_X0Y1_DSP_bot/B3 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ));
 sky130_fd_sc_hd__nand2_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0926_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[3] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0927_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0928_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0929_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0104_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0930_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0072_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0076_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0104_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0066_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ));
 sky130_fd_sc_hd__buf_6 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0931_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0932_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0933_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/A3 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0934_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0935_  (.A(\Tile_X0Y1_DSP_bot/A3 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0110_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0936_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0111_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0937_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0110_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0111_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ));
 sky130_fd_sc_hd__buf_6 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0938_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0939_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ));
 sky130_fd_sc_hd__o2111ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0940_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0941_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0942_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0943_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0118_ ));
 sky130_fd_sc_hd__a22oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0944_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0119_ ));
 sky130_fd_sc_hd__o21bai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0945_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0118_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0119_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ));
 sky130_fd_sc_hd__nand4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0946_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0947_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0120_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0948_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0949_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0950_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0951_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0099_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0952_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0060_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0091_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0090_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0953_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0128_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0954_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0126_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0129_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0955_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0128_ ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0129_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0956_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0131_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0957_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0131_ ),
    .X(\Tile_X0Y1_DSP_bot/Q3 ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0958_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B_N(\Tile_X0Y1_DSP_bot/B3 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0959_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0133_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0960_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0115_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0116_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0105_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0134_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0961_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0133_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0134_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0117_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0962_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0963_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/A4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0964_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0965_  (.A(\Tile_X0Y1_DSP_bot/A4 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0139_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0966_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0140_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0967_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0139_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0140_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ));
 sky130_fd_sc_hd__nor2b_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0968_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B_N(\Tile_X0Y1_DSP_bot/B2 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ));
 sky130_fd_sc_hd__and2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0969_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0970_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0144_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0971_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0144_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0972_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0973_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0974_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0148_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0975_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0109_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0976_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0977_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .B(\Tile_X0Y1_DSP_bot/B4 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0978_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ));
 sky130_fd_sc_hd__a32o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0979_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0980_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0100_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0981_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/B4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ));
 sky130_fd_sc_hd__or4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0982_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0156_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0983_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0156_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ));
 sky130_fd_sc_hd__a221o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0984_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0985_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0148_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0986_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0149_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0114_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0147_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0160_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0987_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0161_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0988_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0145_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0162_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0989_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0161_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0162_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0150_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0990_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0153_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0991_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0160_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0992_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0993_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0994_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0995_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0996_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ));
 sky130_fd_sc_hd__a311o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0997_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0998_  (.A0(\Tile_X0Y1_DSP_bot/C4 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[4] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0172_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_0999_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0172_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1000_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1001_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1002_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0168_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0173_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ));
 sky130_fd_sc_hd__o221a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1003_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0097_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0123_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0124_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0098_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0177_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1004_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0127_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0177_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0125_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1005_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0179_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1006_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0175_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0180_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1007_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0179_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0180_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1008_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0182_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1009_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0182_ ),
    .X(\Tile_X0Y1_DSP_bot/Q4 ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1010_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0178_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0174_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0176_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1011_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0135_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0159_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0165_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ));
 sky130_fd_sc_hd__and4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1012_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0121_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0122_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0167_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0082_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1013_  (.A(\Tile_X0Y1_DSP_bot/A5 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0186_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1014_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1015_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0186_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1016_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1017_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1018_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[0] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1019_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .A2(\Tile_X0Y1_DSP_bot/A5 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0187_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1020_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1021_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0138_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1022_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1023_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/A3 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1024_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1025_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1026_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1027_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1028_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0201_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1029_  (.A(\Tile_X0Y1_DSP_bot/B4 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0202_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1030_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1031_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0202_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1032_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0073_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1033_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1034_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ));
 sky130_fd_sc_hd__or2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1035_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1036_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B5 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1037_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0210_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1038_  (.A(\Tile_X0Y1_DSP_bot/B5 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0211_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1039_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0067_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0212_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1040_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0211_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0212_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1041_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1042_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0028_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1043_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0210_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1044_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0201_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1045_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0190_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0218_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1046_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1047_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0218_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0200_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1048_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1049_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ));
 sky130_fd_sc_hd__o211a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1050_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1051_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1052_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0164_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0163_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0158_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1053_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1054_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1055_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0146_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0198_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1056_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1057_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1058_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ));
 sky130_fd_sc_hd__a41o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1059_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0232_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1060_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0232_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0219_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0233_ ));
 sky130_fd_sc_hd__o41a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1061_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0194_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0234_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1062_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0233_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0234_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1063_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0236_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1064_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0236_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1065_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1066_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1067_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ));
 sky130_fd_sc_hd__o2111ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1068_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0171_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1069_  (.A0(\Tile_X0Y1_DSP_bot/C5 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[5] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0242_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1070_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0242_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ));
 sky130_fd_sc_hd__a21boi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1071_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1072_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0243_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0241_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0240_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1073_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0246_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1074_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0246_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1075_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0248_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1076_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0248_ ),
    .X(\Tile_X0Y1_DSP_bot/Q5 ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1077_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0183_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0245_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0244_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1078_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0224_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0225_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1079_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0221_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0222_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ));
 sky130_fd_sc_hd__a2111o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1080_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0169_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0170_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0252_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1081_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0253_ ));
 sky130_fd_sc_hd__o211ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1082_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0226_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0238_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0254_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1083_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0189_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0229_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1084_  (.A(\Tile_X0Y1_DSP_bot/A6 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0256_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1085_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0024_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1086_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0256_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1087_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1088_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0260_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1089_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0260_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1090_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/A5 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0262_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1091_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0262_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1092_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ));
 sky130_fd_sc_hd__nor2b_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1093_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B_N(\Tile_X0Y1_DSP_bot/A6 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1094_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0266_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1095_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0266_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1096_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0030_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0031_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ));
 sky130_fd_sc_hd__and2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1097_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ));
 sky130_fd_sc_hd__nor2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1098_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .B_N(\Tile_X0Y1_DSP_bot/A4 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1099_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1100_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1101_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .A2(\Tile_X0Y1_DSP_bot/A6 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0257_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1102_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1103_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1104_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1105_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0264_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1106_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0278_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1107_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B2 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0279_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1108_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0278_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0279_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1109_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1110_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1111_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ));
 sky130_fd_sc_hd__a22o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1112_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1113_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ));
 sky130_fd_sc_hd__o2111a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1114_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1115_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0193_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0197_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1116_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0272_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1117_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0277_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0280_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1118_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1119_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1120_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ));
 sky130_fd_sc_hd__or2b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1121_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[6] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ));
 sky130_fd_sc_hd__o21a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1122_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .A2(\Tile_X0Y1_DSP_bot/B6 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1123_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1124_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0040_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0296_ ));
 sky130_fd_sc_hd__a31oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1125_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0206_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0296_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1126_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1127_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B6 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1128_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ));
 sky130_fd_sc_hd__o2bb2a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1129_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1130_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0288_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0302_ ));
 sky130_fd_sc_hd__o22a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1131_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0216_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0220_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1132_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0302_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1133_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1134_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0255_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0276_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0281_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0284_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0285_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ));
 sky130_fd_sc_hd__o211a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1135_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1136_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0227_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0228_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0217_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0308_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1137_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0308_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1138_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1139_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1140_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1141_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1142_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0157_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0237_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0251_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1143_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1144_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0254_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0316_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1145_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1146_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1147_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ));
 sky130_fd_sc_hd__a221oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1148_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0310_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0311_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0317_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0303_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0320_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1149_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0199_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0235_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0306_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0291_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1150_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0312_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0322_ ));
 sky130_fd_sc_hd__o21bai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1151_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0320_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0322_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0314_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0323_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1152_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0323_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0324_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1153_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0252_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0253_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0316_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0324_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1154_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0239_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ));
 sky130_fd_sc_hd__nor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1155_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0298_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0301_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1156_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0304_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0328_ ));
 sky130_fd_sc_hd__a2bb2oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1157_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0328_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1158_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0315_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1159_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0166_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1160_  (.A0(\Tile_X0Y1_DSP_bot/C6 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[6] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0332_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1161_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0332_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1162_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1163_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1164_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0333_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0334_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1165_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0337_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1166_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0337_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0338_ ));
 sky130_fd_sc_hd__xor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1167_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0338_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1168_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0340_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1169_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0340_ ),
    .Y(\Tile_X0Y1_DSP_bot/Q6 ));
 sky130_fd_sc_hd__a32oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1170_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0325_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0336_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0331_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0249_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0335_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1171_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0184_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0185_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0326_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0330_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1172_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B5 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0282_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1173_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0064_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0065_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0344_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1174_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0344_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ));
 sky130_fd_sc_hd__or2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1175_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[7] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0047_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ));
 sky130_fd_sc_hd__o21a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1176_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1177_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1178_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ));
 sky130_fd_sc_hd__and4b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1179_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0350_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1180_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1181_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0049_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0283_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0343_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0352_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1182_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0352_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1183_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0354_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1184_  (.A(\Tile_X0Y1_DSP_bot/A7 ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0355_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1185_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0026_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1186_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0037_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0355_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1187_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0044_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1188_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0191_ ),
    .A2(\Tile_X0Y1_DSP_bot/A7 ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0356_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1189_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1190_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0361_ ));
 sky130_fd_sc_hd__o2111a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1191_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0142_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0143_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1192_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ));
 sky130_fd_sc_hd__o32a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1193_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0268_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0364_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1194_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0361_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0364_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1195_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ));
 sky130_fd_sc_hd__a41o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1196_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0033_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1197_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0032_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1198_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0271_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0363_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1199_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0360_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1200_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1201_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0112_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1202_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B5 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0208_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0373_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1203_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1204_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1205_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0376_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1206_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0373_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0376_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1207_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1208_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1209_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0074_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ));
 sky130_fd_sc_hd__a41o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1210_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ));
 sky130_fd_sc_hd__o22a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1211_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1212_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0375_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ));
 sky130_fd_sc_hd__o2111ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1213_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0384_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1214_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0274_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0259_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1215_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0195_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0287_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0275_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1216_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1217_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0384_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0388_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1218_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1219_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0367_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1220_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1221_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0350_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0354_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0388_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1222_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1223_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1224_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1225_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0378_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0387_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1226_  (.A1(\Tile_X0Y1_DSP_bot/A0 ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0027_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1227_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1228_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1229_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1230_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1231_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0381_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0383_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0402_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1232_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0371_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0403_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1233_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0402_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0403_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0389_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0404_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1234_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0385_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0386_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0290_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0289_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1235_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1236_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0404_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1237_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0397_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0408_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1238_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0408_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0353_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1239_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0321_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ));
 sky130_fd_sc_hd__o32ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1240_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1241_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0412_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1242_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0396_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0406_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0412_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1243_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0400_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0392_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0399_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ));
 sky130_fd_sc_hd__a211oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1244_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0205_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0215_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1245_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1246_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0305_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0329_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ));
 sky130_fd_sc_hd__o221a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1247_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0223_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0250_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0318_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0313_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0418_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1248_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0418_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0419_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1249_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0419_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1250_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1251_  (.A0(\Tile_X0Y1_DSP_bot/C7 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[7] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0422_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1252_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0085_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1253_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0422_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1254_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0425_ ));
 sky130_fd_sc_hd__xor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1255_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0425_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1256_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0427_ ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1257_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0427_ ),
    .X(\Tile_X0Y1_DSP_bot/Q7 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1258_  (.A(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ));
 sky130_fd_sc_hd__or3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1259_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0051_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0297_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ));
 sky130_fd_sc_hd__o311a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1260_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0405_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0393_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0394_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1261_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0286_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0292_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0327_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0309_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1262_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1263_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0433_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1264_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0433_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0434_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1265_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0434_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0416_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0417_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ));
 sky130_fd_sc_hd__o32ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1266_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0431_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0409_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0430_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0429_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0401_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1267_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0395_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0398_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0437_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1268_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1269_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1270_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0070_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1271_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0106_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ));
 sky130_fd_sc_hd__o32ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1272_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0048_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ));
 sky130_fd_sc_hd__o211a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1273_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1274_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1275_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1276_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1277_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0079_ ),
    .B_N(\Tile_X0Y1_DSP_bot/B4 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0447_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1278_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0203_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0447_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1279_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ));
 sky130_fd_sc_hd__nand2_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1280_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1281_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1282_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0141_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ));
 sky130_fd_sc_hd__a32o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1283_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1284_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ));
 sky130_fd_sc_hd__nand2_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1285_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1286_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0440_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0456_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1287_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0368_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0366_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0358_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0456_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1288_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1289_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0369_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0370_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0459_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1290_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0459_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0362_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1291_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ));
 sky130_fd_sc_hd__a22oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1292_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1293_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1294_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1295_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0442_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0444_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0453_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0451_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0465_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1296_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0365_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0377_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0390_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1297_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0465_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1298_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0468_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1299_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0469_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1300_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0374_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0469_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0470_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1301_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B6 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0293_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0471_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1302_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0468_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0470_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0471_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1303_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0380_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0382_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0372_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1304_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1305_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1306_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1307_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0477_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1308_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0041_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1309_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1310_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1311_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1312_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0482_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1313_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0437_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0477_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0482_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1314_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0458_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0460_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1315_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0450_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0446_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0462_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0485_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1316_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0486_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1317_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0485_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0486_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ));
 sky130_fd_sc_hd__a21o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1318_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1319_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0474_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0475_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0489_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1320_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0391_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0407_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0489_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ));
 sky130_fd_sc_hd__a31o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1321_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0029_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0349_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0345_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ));
 sky130_fd_sc_hd__a21o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1322_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1323_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1324_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ));
 sky130_fd_sc_hd__a221o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1325_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0432_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1326_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1327_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0495_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1328_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1329_  (.A0(\Tile_X0Y1_DSP_bot/C8 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[8] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0499_ ));
 sky130_fd_sc_hd__or2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1330_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ),
    .B_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0500_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1331_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0499_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0500_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1332_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ));
 sky130_fd_sc_hd__or3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1333_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0503_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1334_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0503_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1335_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0307_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0413_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0415_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1336_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0410_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0411_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0506_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1337_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0319_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0506_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0342_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0507_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1338_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0420_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0507_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1339_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0421_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0424_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1340_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1341_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1342_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0510_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0504_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1343_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0513_ ));
 sky130_fd_sc_hd__a31o_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1344_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0513_ ),
    .X(\Tile_X0Y1_DSP_bot/Q8 ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1345_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0341_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0508_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0509_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0514_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1346_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0501_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0497_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0496_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0515_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1347_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0514_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0502_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0515_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ));
 sky130_fd_sc_hd__a32oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1348_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0505_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0414_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0517_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1349_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0436_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0518_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1350_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0517_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0492_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0518_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1351_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ));
 sky130_fd_sc_hd__buf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1352_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1353_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1354_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0188_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ));
 sky130_fd_sc_hd__nand4_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1355_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1356_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .A2(\Tile_X0Y1_DSP_bot/A4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0213_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1357_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1358_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0102_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0204_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1359_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1360_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1361_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0524_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1362_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1363_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0071_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0441_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0532_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1364_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0532_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ));
 sky130_fd_sc_hd__a221oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1365_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ));
 sky130_fd_sc_hd__o22a_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1366_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0522_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0526_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0528_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1367_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ));
 sky130_fd_sc_hd__a211o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1368_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0045_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0537_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1369_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0530_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0531_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0538_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1370_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0537_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0538_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1371_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0540_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1372_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0448_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0541_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1373_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0107_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0196_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0542_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1374_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0540_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0541_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0542_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1375_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0449_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0544_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1376_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0299_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0445_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0544_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0452_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1377_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0546_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1378_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0547_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1379_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0546_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0547_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0548_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1380_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0548_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1381_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0550_ ));
 sky130_fd_sc_hd__a21oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1382_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0455_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0454_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0550_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ));
 sky130_fd_sc_hd__o2bb2a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1383_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0063_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1384_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0207_ ),
    .A2(\Tile_X0Y1_DSP_bot/B7 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0075_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0346_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1385_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ));
 sky130_fd_sc_hd__nor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1386_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1387_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1388_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1389_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0487_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0466_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0476_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ));
 sky130_fd_sc_hd__a221o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1390_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0463_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0457_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0529_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0443_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1391_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0555_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ));
 sky130_fd_sc_hd__o22ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1392_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0551_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0534_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1393_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1394_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0478_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0473_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0472_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1395_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1396_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0565_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1397_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0493_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0565_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1398_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0479_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0480_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0567_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1399_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0567_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0467_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0481_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0464_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0568_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1400_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0568_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ));
 sky130_fd_sc_hd__o211a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1401_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0484_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0558_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0560_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0561_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1402_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0571_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1403_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0483_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0491_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0490_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1404_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0571_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1405_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1406_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1407_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0520_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0574_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1408_  (.A0(\Tile_X0Y1_DSP_bot/C9 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[9] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0577_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1409_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0577_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ));
 sky130_fd_sc_hd__o21bai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1410_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1411_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0575_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0576_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0580_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1412_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0580_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0578_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1413_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0582_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1414_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0583_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1415_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0582_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0583_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1416_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0585_ ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1417_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0585_ ),
    .X(\Tile_X0Y1_DSP_bot/Q9 ));
 sky130_fd_sc_hd__o21a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1418_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0564_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0566_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1419_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0587_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1420_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0588_ ));
 sky130_fd_sc_hd__nand3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1421_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0557_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0589_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1422_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0588_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0589_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0590_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1423_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0572_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0590_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0494_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1424_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0592_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1425_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0593_ ));
 sky130_fd_sc_hd__a221o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1426_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0230_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0593_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1427_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0525_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0523_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0527_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0595_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1428_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .A2(\Tile_X0Y1_DSP_bot/A4 ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0136_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0595_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1429_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1430_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0113_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1431_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0258_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0357_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1432_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0359_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1433_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0601_ ));
 sky130_fd_sc_hd__o2111ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1434_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0600_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0602_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1435_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0601_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0602_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1436_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ));
 sky130_fd_sc_hd__or4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1437_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0050_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0080_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1438_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0606_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1439_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0606_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1440_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0439_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0608_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1441_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0605_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0533_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0603_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1442_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0608_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1443_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ));
 sky130_fd_sc_hd__nand3_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1444_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ));
 sky130_fd_sc_hd__a21boi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1445_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0553_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0545_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0543_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ));
 sky130_fd_sc_hd__a21boi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1446_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1447_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0552_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0554_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0535_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0539_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0559_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0615_ ));
 sky130_fd_sc_hd__a41oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1448_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0461_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0488_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0556_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0615_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ));
 sky130_fd_sc_hd__nand3b_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1449_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1450_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1451_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0607_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0610_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0549_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ));
 sky130_fd_sc_hd__nor3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1452_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ),
    .C_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0620_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1453_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0563_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0569_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0562_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0621_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1454_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0620_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0621_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ));
 sky130_fd_sc_hd__o21ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1455_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ));
 sky130_fd_sc_hd__a21o_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1456_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0587_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0592_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ));
 sky130_fd_sc_hd__a32oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1457_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1458_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1459_  (.A0(\Tile_X0Y1_DSP_bot/C10 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[10] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0086_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0627_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1460_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0627_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1461_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1462_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1463_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0628_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0629_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1464_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1465_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1466_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1467_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0635_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1468_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0630_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0635_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0579_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1469_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0637_ ));
 sky130_fd_sc_hd__a31o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1470_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0637_ ),
    .X(\Tile_X0Y1_DSP_bot/Q10 ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1471_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0624_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0626_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0631_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1472_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0516_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0581_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0633_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1473_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0611_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0640_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1474_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0570_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0616_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0617_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0640_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1475_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0642_ ));
 sky130_fd_sc_hd__a31o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1476_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0643_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1477_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0209_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1478_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0155_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1479_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0265_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0267_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1480_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/A7 ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0647_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1481_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0025_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0648_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1482_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0101_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0132_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0647_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0648_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1483_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1484_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ));
 sky130_fd_sc_hd__o211ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1485_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0192_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0599_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ));
 sky130_fd_sc_hd__and4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1486_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0103_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0653_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1487_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0649_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0650_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0654_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1488_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0261_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0263_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ));
 sky130_fd_sc_hd__o21bai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1489_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0653_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0654_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ));
 sky130_fd_sc_hd__o2111ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1490_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0269_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0270_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0347_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1491_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0652_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ));
 sky130_fd_sc_hd__o211ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1492_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0659_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1493_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0379_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0214_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ));
 sky130_fd_sc_hd__a32o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1494_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0151_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0152_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1495_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0662_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1496_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0643_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0659_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0662_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1497_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0644_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0645_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1498_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0657_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0658_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0661_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ));
 sky130_fd_sc_hd__a31oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1499_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0597_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0598_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0604_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0609_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1500_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1501_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0594_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0668_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1502_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0108_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0668_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0596_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ));
 sky130_fd_sc_hd__a21boi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1503_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1504_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0613_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0619_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0612_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ));
 sky130_fd_sc_hd__nand3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1505_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1506_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1507_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0667_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1508_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1509_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1510_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0642_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1511_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0676_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0678_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1512_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0614_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0618_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0623_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0625_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0678_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1513_  (.A0(\Tile_X0Y1_DSP_bot/C11 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[11] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0680_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1514_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1515_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0680_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1516_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1517_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ));
 sky130_fd_sc_hd__nor4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1518_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0685_ ));
 sky130_fd_sc_hd__o22a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1519_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0638_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0684_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0686_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1520_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0685_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0686_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1521_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0688_ ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1522_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0688_ ),
    .X(\Tile_X0Y1_DSP_bot/Q11 ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1523_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0677_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0679_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0682_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ));
 sky130_fd_sc_hd__a31oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1524_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ));
 sky130_fd_sc_hd__o2111a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1525_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0675_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0622_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1526_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0435_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0519_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0586_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1527_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0674_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0672_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0671_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0693_ ));
 sky130_fd_sc_hd__o22ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1528_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0670_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0673_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0693_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0641_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0694_ ));
 sky130_fd_sc_hd__a31oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1529_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0691_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0591_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0573_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0694_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ));
 sky130_fd_sc_hd__or2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1530_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1531_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1532_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1533_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1534_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ));
 sky130_fd_sc_hd__nand4_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1535_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0295_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0698_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ));
 sky130_fd_sc_hd__and3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1536_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1537_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0700_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ));
 sky130_fd_sc_hd__o311a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1538_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0154_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0646_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0655_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0651_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0704_ ));
 sky130_fd_sc_hd__o31a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1539_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0137_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0704_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0656_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1540_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ));
 sky130_fd_sc_hd__nor3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1541_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0705_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0703_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1542_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0664_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0665_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0666_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0708_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1543_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0669_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0708_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0663_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1544_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0710_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1545_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0709_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0706_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1546_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1547_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0710_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1548_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1549_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1550_  (.A0(\Tile_X0Y1_DSP_bot/C12 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[12] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0716_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1551_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0716_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1552_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1553_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1554_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1555_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0715_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0719_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1556_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1557_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1558_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0724_ ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1559_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0724_ ),
    .X(\Tile_X0Y1_DSP_bot/Q12 ));
 sky130_fd_sc_hd__a21oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1560_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1561_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0726_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1562_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0727_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1563_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0521_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0726_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0727_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ));
 sky130_fd_sc_hd__xor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1564_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1565_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0696_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0699_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1566_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0660_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0731_ ));
 sky130_fd_sc_hd__a311o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1567_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0231_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0697_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0348_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0731_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0729_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ));
 sky130_fd_sc_hd__a211oi_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1568_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ));
 sky130_fd_sc_hd__o211a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1569_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0702_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0707_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0732_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1570_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0735_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1571_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0735_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1572_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0712_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0714_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1573_  (.A0(\Tile_X0Y1_DSP_bot/C13 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[13] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0738_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1574_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0738_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1575_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1576_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1577_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0739_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0740_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0742_ ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1578_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0736_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0737_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0742_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1579_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ));
 sky130_fd_sc_hd__a21bo_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1580_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0690_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0721_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0720_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0745_ ));
 sky130_fd_sc_hd__xor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1581_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0745_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1582_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ),
    .S(\Tile_X0Y1_DSP_bot/ConfigBits[5] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0747_ ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1583_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0747_ ),
    .X(\Tile_X0Y1_DSP_bot/Q13 ));
 sky130_fd_sc_hd__a211o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1584_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0536_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0294_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1585_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1586_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1587_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0748_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0749_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1588_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0711_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1589_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0753_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1590_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0754_ ));
 sky130_fd_sc_hd__o221ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1591_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0753_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0754_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1592_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0756_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1593_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0734_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0757_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1594_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0756_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0757_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0758_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1595_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0750_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0751_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0759_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1596_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0733_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0752_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0758_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0759_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1597_  (.A0(\Tile_X0Y1_DSP_bot/C14 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[14] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0761_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1598_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0761_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1599_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1600_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1601_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1602_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0713_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0692_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0695_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0766_ ));
 sky130_fd_sc_hd__o41ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1603_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0725_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0766_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0717_ ),
    .A4(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0718_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0743_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1604_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0632_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0689_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0768_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1605_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0722_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0683_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0769_ ));
 sky130_fd_sc_hd__o211ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1606_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0768_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0639_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0769_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0744_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ));
 sky130_fd_sc_hd__a21boi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1607_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1608_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0772_ ));
 sky130_fd_sc_hd__and2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1609_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ));
 sky130_fd_sc_hd__a2bb2o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1610_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0772_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .X(\Tile_X0Y1_DSP_bot/Q14 ));
 sky130_fd_sc_hd__o221a_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1611_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0273_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0300_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0701_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0728_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0730_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ));
 sky130_fd_sc_hd__o31ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1612_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1613_  (.A0(\Tile_X0Y1_DSP_bot/C15 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[15] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0776_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1614_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0776_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0423_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1615_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1616_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0779_ ));
 sky130_fd_sc_hd__o311ai_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1617_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0351_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0438_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0774_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0779_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ));
 sky130_fd_sc_hd__o2111a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1618_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .D1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0781_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1619_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0782_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1620_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0765_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0771_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1621_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0782_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0784_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1622_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0781_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0784_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1623_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0786_ ));
 sky130_fd_sc_hd__o21ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1624_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0786_ ),
    .Y(\Tile_X0Y1_DSP_bot/Q15 ));
 sky130_fd_sc_hd__nand2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1625_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1626_  (.A0(\Tile_X0Y1_DSP_bot/C16 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[16] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0788_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1627_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0788_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ));
 sky130_fd_sc_hd__xnor2_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1628_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1629_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0741_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0767_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0791_ ));
 sky130_fd_sc_hd__a32oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1630_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0755_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0760_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0762_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0777_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0792_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1631_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0791_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0792_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0793_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1632_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0763_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0764_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0778_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0794_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1633_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0780_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0793_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0794_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0770_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1634_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1635_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0797_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1636_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0797_ ),
    .X(\Tile_X0Y1_DSP_bot/Q16 ));
 sky130_fd_sc_hd__nand3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1637_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0789_ ),
    .C(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ));
 sky130_fd_sc_hd__nand2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1638_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1639_  (.A0(\Tile_X0Y1_DSP_bot/C17 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[17] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0800_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1640_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0800_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ));
 sky130_fd_sc_hd__a221o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1641_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B2(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1642_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0801_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1643_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ));
 sky130_fd_sc_hd__a22o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1644_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ));
 sky130_fd_sc_hd__nand4_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1645_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0804_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1646_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0807_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1647_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0807_ ),
    .X(\Tile_X0Y1_DSP_bot/Q17 ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1648_  (.A0(\Tile_X0Y1_DSP_bot/C18 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[18] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0808_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1649_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0808_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1650_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1651_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .A2(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0811_ ));
 sky130_fd_sc_hd__or2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1652_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0812_ ));
 sky130_fd_sc_hd__nand3_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1653_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0795_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0790_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0802_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ));
 sky130_fd_sc_hd__o21a_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1654_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0803_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0798_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ));
 sky130_fd_sc_hd__a22oi_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1655_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0811_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0812_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1656_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .A2(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1657_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .C(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1658_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ));
 sky130_fd_sc_hd__a31o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1659_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .A3(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0819_ ));
 sky130_fd_sc_hd__a2bb2o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1660_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0819_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0021_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ),
    .X(\Tile_X0Y1_DSP_bot/Q18 ));
 sky130_fd_sc_hd__inv_2 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1661_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0820_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1662_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0775_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0809_ ),
    .C(\Tile_X0Y1_DSP_bot/ConfigBits[4] ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0821_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1663_  (.A0(\Tile_X0Y1_DSP_bot/C19 ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[19] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0498_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0822_ ));
 sky130_fd_sc_hd__mux2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1664_  (.A0(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0822_ ),
    .A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ),
    .S(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0681_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0823_ ));
 sky130_fd_sc_hd__xnor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1665_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0823_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ));
 sky130_fd_sc_hd__o21bai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1666_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0821_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ),
    .B1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1667_  (.A1_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .A2_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0817_ ),
    .B2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0816_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0826_ ));
 sky130_fd_sc_hd__o211ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1668_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0787_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0810_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0824_ ),
    .C1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0826_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ));
 sky130_fd_sc_hd__a21o_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1669_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0094_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0828_ ));
 sky130_fd_sc_hd__o21ai_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1670_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0428_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0820_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0828_ ),
    .Y(\Tile_X0Y1_DSP_bot/Q19 ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1671_  (.A(\Tile_X0Y1_DSP_bot/clr ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1672_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0034_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0035_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0000_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1673_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0058_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0001_ ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1674_  (.A(\Tile_X0Y1_DSP_bot/clr ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1675_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0093_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0831_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1676_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0831_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0002_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1677_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0130_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0832_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1678_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0832_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0003_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1679_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0181_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0833_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1680_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0833_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0004_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1681_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0247_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0834_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1682_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0834_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0005_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1683_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0339_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0006_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1684_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0426_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0835_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1685_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0835_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0007_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1686_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0511_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0512_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0836_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1687_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0836_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0008_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1688_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0584_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0837_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1689_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0837_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0009_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1690_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0634_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0636_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0838_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1691_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0838_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0010_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1692_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0687_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0839_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1693_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0839_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0011_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1694_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0723_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0840_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1695_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0840_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0012_ ));
 sky130_fd_sc_hd__and2b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1696_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0746_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0841_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1697_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0841_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0013_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1698_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0783_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0773_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0014_ ));
 sky130_fd_sc_hd__nor2_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1699_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0785_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0015_ ));
 sky130_fd_sc_hd__and3b_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1700_  (.A_N(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0830_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0799_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0796_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0842_ ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1701_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0842_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0016_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1702_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0805_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0806_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0017_ ));
 sky130_fd_sc_hd__and3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1703_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0813_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0814_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0818_ ),
    .X(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0020_ ));
 sky130_fd_sc_hd__nor3_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1704_  (.A(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .B(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0020_ ),
    .C(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0815_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0018_ ));
 sky130_fd_sc_hd__a21oi_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1705_  (.A1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0825_ ),
    .A2(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0827_ ),
    .B1(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0829_ ),
    .Y(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0019_ ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1706_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0000_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1707_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0001_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1708_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0002_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1709_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0003_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1710_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0004_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1711_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0005_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1712_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0006_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1713_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0007_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1714_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0008_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[8] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1715_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0009_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[9] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1716_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0010_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[10] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1717_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0011_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[11] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1718_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0012_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[12] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1719_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0013_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[13] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1720_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0014_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[14] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1721_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0015_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[15] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1722_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0016_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[16] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1723_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0017_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[17] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1724_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0018_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[18] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1725_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/Inst_MULADD/_0019_ ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/ACC[19] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1726_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A0 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1727_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A1 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1728_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A2 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1729_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A3 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1730_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A4 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1731_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A5 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1732_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A6 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1733_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/A7 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/A_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1734_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B0 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1735_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B1 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1736_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B2 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1737_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B3 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1738_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B4 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1739_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B5 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1740_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B6 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1741_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/B7 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/B_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1742_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C0 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1743_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C1 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1744_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C2 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1745_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C3 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1746_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C4 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1747_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C5 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1748_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C6 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1749_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C7 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1750_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C8 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1751_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C9 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1752_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C10 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1753_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C11 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1754_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C12 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1755_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C13 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1756_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C14 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1757_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C15 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1758_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C16 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1759_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C17 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1760_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C18 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 \Tile_X0Y1_DSP_bot/Inst_MULADD/_1761_  (.CLK(net333),
    .D(\Tile_X0Y1_DSP_bot/C19 ),
    .Q(\Tile_X0Y1_DSP_bot/Inst_MULADD/C_reg[19] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[0] ),
    .X(\Tile_X0Y1_N4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[1] ),
    .X(\Tile_X0Y1_N4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[10] ),
    .X(\Tile_X0Y1_N4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[11] ),
    .X(\Tile_X0Y1_N4BEG[11] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[2] ),
    .X(\Tile_X0Y1_N4BEG[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[3] ),
    .X(\Tile_X0Y1_N4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[4] ),
    .X(\Tile_X0Y1_N4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[5] ),
    .X(\Tile_X0Y1_N4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[6] ),
    .X(\Tile_X0Y1_N4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[7] ),
    .X(\Tile_X0Y1_N4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[8] ),
    .X(\Tile_X0Y1_N4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/N4BEG_i[9] ),
    .X(\Tile_X0Y1_N4BEG[9] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/N4END_inbuf_0/_0_  (.A(net311),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_1/_0_  (.A(net312),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_10/_0_  (.A(net306),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[10] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_11/_0_  (.A(net307),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_2/_0_  (.A(net313),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/N4END_inbuf_3/_0_  (.A(net314),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_4/_0_  (.A(net315),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_5/_0_  (.A(net316),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[5] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_6/_0_  (.A(net302),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_7/_0_  (.A(net303),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_8/_0_  (.A(net304),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/N4END_inbuf_9/_0_  (.A(net305),
    .X(\Tile_X0Y1_DSP_bot/N4BEG_i[9] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[0] ),
    .X(\Tile_X0Y1_NN4BEG[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[1] ),
    .X(\Tile_X0Y1_NN4BEG[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[10] ),
    .X(\Tile_X0Y1_NN4BEG[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[11] ),
    .X(\Tile_X0Y1_NN4BEG[11] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[2] ),
    .X(\Tile_X0Y1_NN4BEG[2] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[3] ),
    .X(\Tile_X0Y1_NN4BEG[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[4] ),
    .X(\Tile_X0Y1_NN4BEG[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[5] ),
    .X(\Tile_X0Y1_NN4BEG[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[6] ),
    .X(\Tile_X0Y1_NN4BEG[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[7] ),
    .X(\Tile_X0Y1_NN4BEG[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[8] ),
    .X(\Tile_X0Y1_NN4BEG[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/NN4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/NN4BEG_i[9] ),
    .X(\Tile_X0Y1_NN4BEG[9] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/NN4END_inbuf_0/_0_  (.A(net327),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_1/_0_  (.A(net328),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_10/_0_  (.A(net322),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_11/_0_  (.A(net323),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_2/_0_  (.A(net329),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[2] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_3/_0_  (.A(net330),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_4/_0_  (.A(net331),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_5/_0_  (.A(net332),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_6/_0_  (.A(net318),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_7/_0_  (.A(net319),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_8/_0_  (.A(net320),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/NN4END_inbuf_9/_0_  (.A(net321),
    .X(\Tile_X0Y1_DSP_bot/NN4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[0] ),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[1] ),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[11] ),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[2] ),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[3] ),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[4] ),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[5] ),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[6] ),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[7] ),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[8] ),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/S4BEG_i[9] ),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/S4END_inbuf_0/_0_  (.A(\Tile_X0Y0_S4BEG[4] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_1/_0_  (.A(\Tile_X0Y0_S4BEG[5] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_10/_0_  (.A(\Tile_X0Y0_S4BEG[14] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_11/_0_  (.A(\Tile_X0Y0_S4BEG[15] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4END_inbuf_2/_0_  (.A(\Tile_X0Y0_S4BEG[6] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_3/_0_  (.A(\Tile_X0Y0_S4BEG[7] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_4/_0_  (.A(\Tile_X0Y0_S4BEG[8] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[4] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/S4END_inbuf_5/_0_  (.A(\Tile_X0Y0_S4BEG[9] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[5] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/S4END_inbuf_6/_0_  (.A(\Tile_X0Y0_S4BEG[10] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/S4END_inbuf_7/_0_  (.A(\Tile_X0Y0_S4BEG[11] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_8/_0_  (.A(\Tile_X0Y0_S4BEG[12] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[8] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/S4END_inbuf_9/_0_  (.A(\Tile_X0Y0_S4BEG[13] ),
    .X(\Tile_X0Y1_DSP_bot/S4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[0] ),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[1] ),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[10] ),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[11] ),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[2] ),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[3] ),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[4] ),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[5] ),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[6] ),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[7] ),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[8] ),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/SS4BEG_i[9] ),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_0/_0_  (.A(\Tile_X0Y0_SS4BEG[4] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_1/_0_  (.A(\Tile_X0Y0_SS4BEG[5] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/SS4END_inbuf_10/_0_  (.A(\Tile_X0Y0_SS4BEG[14] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/SS4END_inbuf_11/_0_  (.A(\Tile_X0Y0_SS4BEG[15] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_2/_0_  (.A(\Tile_X0Y0_SS4BEG[6] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_3/_0_  (.A(\Tile_X0Y0_SS4BEG[7] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_4/_0_  (.A(\Tile_X0Y0_SS4BEG[8] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_5/_0_  (.A(\Tile_X0Y0_SS4BEG[9] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_6/_0_  (.A(\Tile_X0Y0_SS4BEG[10] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/SS4END_inbuf_7/_0_  (.A(\Tile_X0Y0_SS4BEG[11] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[7] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/SS4END_inbuf_8/_0_  (.A(\Tile_X0Y0_SS4BEG[12] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/SS4END_inbuf_9/_0_  (.A(\Tile_X0Y0_SS4BEG[13] ),
    .X(\Tile_X0Y1_DSP_bot/SS4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[0] ),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[1] ),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[2] ),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[3] ),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[4] ),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[5] ),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[6] ),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[7] ),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[8] ),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/W6BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/W6BEG_i[9] ),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_0/_0_  (.A(net358),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_1/_0_  (.A(net359),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_2/_0_  (.A(net360),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_3/_0_  (.A(net361),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_4/_0_  (.A(net362),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_5/_0_  (.A(net363),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_6/_0_  (.A(net364),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_7/_0_  (.A(net365),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_8/_0_  (.A(net355),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/W6END_inbuf_9/_0_  (.A(net356),
    .X(\Tile_X0Y1_DSP_bot/W6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[0] ),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[1] ),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[10] ),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[11] ),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[2] ),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[3] ),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[4] ),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[5] ),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[6] ),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[7] ),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[8] ),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/WW4BEG_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/WW4BEG_i[9] ),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_0/_0_  (.A(net376),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_1/_0_  (.A(net377),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_10/_0_  (.A(net371),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_11/_0_  (.A(net372),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_2/_0_  (.A(net378),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_3/_0_  (.A(net379),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_4/_0_  (.A(net380),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_5/_0_  (.A(net381),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_6/_0_  (.A(net367),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_7/_0_  (.A(net368),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_8/_0_  (.A(net369),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/WW4END_inbuf_9/_0_  (.A(net370),
    .X(\Tile_X0Y1_DSP_bot/WW4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_0/_0_  (.A(net229),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_1/_0_  (.A(net240),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_10/_0_  (.A(net230),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_11/_0_  (.A(net231),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_12/_0_  (.A(net232),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[12] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/data_inbuf_13/_0_  (.A(net233),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_14/_0_  (.A(net234),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_15/_0_  (.A(net235),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_16/_0_  (.A(net236),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_17/_0_  (.A(net237),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_18/_0_  (.A(net238),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_19/_0_  (.A(net239),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_2/_0_  (.A(net251),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_20/_0_  (.A(net241),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[20] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_21/_0_  (.A(net242),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_22/_0_  (.A(net243),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_23/_0_  (.A(net244),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_24/_0_  (.A(net245),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_25/_0_  (.A(net246),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_26/_0_  (.A(net247),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_27/_0_  (.A(net248),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_28/_0_  (.A(net249),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_29/_0_  (.A(net250),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_3/_0_  (.A(net254),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_30/_0_  (.A(net252),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[30] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_31/_0_  (.A(net253),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_4/_0_  (.A(net255),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_5/_0_  (.A(net256),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_6/_0_  (.A(net257),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_7/_0_  (.A(net258),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_8/_0_  (.A(net259),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_inbuf_9/_0_  (.A(net260),
    .X(\Tile_X0Y1_DSP_bot/FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[0] ),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[1] ),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[10] ),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[11] ),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_12/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[12] ),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_13/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[13] ),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_14/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[14] ),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_15/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[15] ),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_16/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[16] ),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_17/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[17] ),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_18/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[18] ),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_19/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[19] ),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[2] ),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_20/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[20] ),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_21/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[21] ),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_22/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[22] ),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_23/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[23] ),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_24/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[24] ),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_25/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[25] ),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_26/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[26] ),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_27/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[27] ),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_28/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[28] ),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_29/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[29] ),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[3] ),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_30/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[30] ),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_31/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[31] ),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[4] ),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[5] ),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[6] ),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[7] ),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[8] ),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/data_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameData_O_i[9] ),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/inst_clk_buf  (.A(net333),
    .X(Tile_X0Y1_UserCLKo));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_0/_0_  (.A(net261),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_1/_0_  (.A(net272),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_10/_0_  (.A(net262),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_11/_0_  (.A(net263),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_12/_0_  (.A(net264),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_13/_0_  (.A(net265),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_14/_0_  (.A(net266),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_15/_0_  (.A(net267),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_16/_0_  (.A(net268),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_17/_0_  (.A(net269),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_18/_0_  (.A(net270),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_19/_0_  (.A(net271),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_2/_0_  (.A(net273),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_3/_0_  (.A(net274),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_4/_0_  (.A(net275),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_5/_0_  (.A(net276),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_6/_0_  (.A(net277),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_7/_0_  (.A(net278),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__buf_1 \Tile_X0Y1_DSP_bot/strobe_inbuf_8/_0_  (.A(net279),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \Tile_X0Y1_DSP_bot/strobe_inbuf_9/_0_  (.A(net280),
    .X(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_0/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[0] ),
    .X(\Tile_X0Y1_FrameStrobe_O[0] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_1/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[1] ),
    .X(\Tile_X0Y1_FrameStrobe_O[1] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_10/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[10] ),
    .X(\Tile_X0Y1_FrameStrobe_O[10] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_11/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[11] ),
    .X(\Tile_X0Y1_FrameStrobe_O[11] ));
 sky130_fd_sc_hd__clkbuf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_12/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[12] ),
    .X(\Tile_X0Y1_FrameStrobe_O[12] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_13/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[13] ),
    .X(\Tile_X0Y1_FrameStrobe_O[13] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_14/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[14] ),
    .X(\Tile_X0Y1_FrameStrobe_O[14] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_15/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[15] ),
    .X(\Tile_X0Y1_FrameStrobe_O[15] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/strobe_outbuf_16/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[16] ),
    .X(\Tile_X0Y1_FrameStrobe_O[16] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_17/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[17] ),
    .X(\Tile_X0Y1_FrameStrobe_O[17] ));
 sky130_fd_sc_hd__buf_2 \Tile_X0Y1_DSP_bot/strobe_outbuf_18/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[18] ),
    .X(\Tile_X0Y1_FrameStrobe_O[18] ));
 sky130_fd_sc_hd__clkbuf_4 \Tile_X0Y1_DSP_bot/strobe_outbuf_19/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[19] ),
    .X(\Tile_X0Y1_FrameStrobe_O[19] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_2/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[2] ),
    .X(\Tile_X0Y1_FrameStrobe_O[2] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_3/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[3] ),
    .X(\Tile_X0Y1_FrameStrobe_O[3] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_4/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[4] ),
    .X(\Tile_X0Y1_FrameStrobe_O[4] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_5/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[5] ),
    .X(\Tile_X0Y1_FrameStrobe_O[5] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_6/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[6] ),
    .X(\Tile_X0Y1_FrameStrobe_O[6] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_7/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[7] ),
    .X(\Tile_X0Y1_FrameStrobe_O[7] ));
 sky130_fd_sc_hd__buf_12 \Tile_X0Y1_DSP_bot/strobe_outbuf_8/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[8] ),
    .X(\Tile_X0Y1_FrameStrobe_O[8] ));
 sky130_fd_sc_hd__buf_8 \Tile_X0Y1_DSP_bot/strobe_outbuf_9/_0_  (.A(\Tile_X0Y1_DSP_bot/FrameStrobe_O_i[9] ),
    .X(\Tile_X0Y1_FrameStrobe_O[9] ));
 sky130_fd_sc_hd__buf_4 input1 (.A(Tile_X0Y0_E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(Tile_X0Y0_E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(Tile_X0Y0_S2MID[7]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(Tile_X0Y0_S4END[0]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(Tile_X0Y0_S4END[10]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(Tile_X0Y0_S4END[11]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(Tile_X0Y0_S4END[12]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(Tile_X0Y0_S4END[13]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(Tile_X0Y0_S4END[14]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(Tile_X0Y0_S4END[15]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(Tile_X0Y0_S4END[1]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(Tile_X0Y0_S4END[2]),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(Tile_X0Y0_E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(Tile_X0Y0_S4END[3]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(Tile_X0Y0_S4END[4]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(Tile_X0Y0_S4END[5]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(Tile_X0Y0_S4END[6]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(Tile_X0Y0_S4END[7]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(Tile_X0Y0_S4END[8]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(Tile_X0Y0_S4END[9]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(Tile_X0Y0_SS4END[0]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(Tile_X0Y0_SS4END[10]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(Tile_X0Y0_SS4END[11]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(Tile_X0Y0_E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(Tile_X0Y0_SS4END[12]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(Tile_X0Y0_SS4END[13]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(Tile_X0Y0_SS4END[14]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(Tile_X0Y0_SS4END[15]),
    .X(net123));
 sky130_fd_sc_hd__buf_2 input124 (.A(Tile_X0Y0_SS4END[1]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(Tile_X0Y0_SS4END[2]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(Tile_X0Y0_SS4END[3]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(Tile_X0Y0_SS4END[4]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(Tile_X0Y0_SS4END[5]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(Tile_X0Y0_SS4END[6]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input13 (.A(Tile_X0Y0_E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(Tile_X0Y0_SS4END[7]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(Tile_X0Y0_SS4END[8]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(Tile_X0Y0_SS4END[9]),
    .X(net132));
 sky130_fd_sc_hd__buf_4 input133 (.A(Tile_X0Y0_W1END[0]),
    .X(net133));
 sky130_fd_sc_hd__buf_4 input134 (.A(Tile_X0Y0_W1END[1]),
    .X(net134));
 sky130_fd_sc_hd__buf_4 input135 (.A(Tile_X0Y0_W1END[2]),
    .X(net135));
 sky130_fd_sc_hd__buf_4 input136 (.A(Tile_X0Y0_W1END[3]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(Tile_X0Y0_W2END[0]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(Tile_X0Y0_W2END[1]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(Tile_X0Y0_W2END[2]),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(Tile_X0Y0_E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input140 (.A(Tile_X0Y0_W2END[3]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(Tile_X0Y0_W2END[4]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(Tile_X0Y0_W2END[5]),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 input143 (.A(Tile_X0Y0_W2END[6]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 input144 (.A(Tile_X0Y0_W2END[7]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(Tile_X0Y0_W2MID[0]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(Tile_X0Y0_W2MID[1]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 input147 (.A(Tile_X0Y0_W2MID[2]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 input148 (.A(Tile_X0Y0_W2MID[3]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(Tile_X0Y0_W2MID[4]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(Tile_X0Y0_E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input150 (.A(Tile_X0Y0_W2MID[5]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 input151 (.A(Tile_X0Y0_W2MID[6]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(Tile_X0Y0_W2MID[7]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(Tile_X0Y0_W6END[0]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(Tile_X0Y0_W6END[10]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(Tile_X0Y0_W6END[11]),
    .X(net155));
 sky130_fd_sc_hd__buf_4 input156 (.A(Tile_X0Y0_W6END[1]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 input157 (.A(Tile_X0Y0_W6END[2]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(Tile_X0Y0_W6END[3]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(Tile_X0Y0_W6END[4]),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input16 (.A(Tile_X0Y0_E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(Tile_X0Y0_W6END[5]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(Tile_X0Y0_W6END[6]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(Tile_X0Y0_W6END[7]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(Tile_X0Y0_W6END[8]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(Tile_X0Y0_W6END[9]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(Tile_X0Y0_WW4END[0]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(Tile_X0Y0_WW4END[10]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(Tile_X0Y0_WW4END[11]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(Tile_X0Y0_WW4END[12]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(Tile_X0Y0_WW4END[13]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(Tile_X0Y0_E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(Tile_X0Y0_WW4END[14]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(Tile_X0Y0_WW4END[15]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(Tile_X0Y0_WW4END[1]),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(Tile_X0Y0_WW4END[2]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(Tile_X0Y0_WW4END[3]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(Tile_X0Y0_WW4END[4]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(Tile_X0Y0_WW4END[5]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(Tile_X0Y0_WW4END[6]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(Tile_X0Y0_WW4END[7]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(Tile_X0Y0_WW4END[8]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(Tile_X0Y0_E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(Tile_X0Y0_WW4END[9]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(Tile_X0Y1_E1END[0]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 input182 (.A(Tile_X0Y1_E1END[1]),
    .X(net182));
 sky130_fd_sc_hd__buf_4 input183 (.A(Tile_X0Y1_E1END[2]),
    .X(net183));
 sky130_fd_sc_hd__buf_4 input184 (.A(Tile_X0Y1_E1END[3]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(Tile_X0Y1_E2END[0]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(Tile_X0Y1_E2END[1]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 input187 (.A(Tile_X0Y1_E2END[2]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 input188 (.A(Tile_X0Y1_E2END[3]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 input189 (.A(Tile_X0Y1_E2END[4]),
    .X(net189));
 sky130_fd_sc_hd__buf_2 input19 (.A(Tile_X0Y0_E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(Tile_X0Y1_E2END[5]),
    .X(net190));
 sky130_fd_sc_hd__buf_2 input191 (.A(Tile_X0Y1_E2END[6]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(Tile_X0Y1_E2END[7]),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input193 (.A(Tile_X0Y1_E2MID[0]),
    .X(net193));
 sky130_fd_sc_hd__buf_2 input194 (.A(Tile_X0Y1_E2MID[1]),
    .X(net194));
 sky130_fd_sc_hd__buf_2 input195 (.A(Tile_X0Y1_E2MID[2]),
    .X(net195));
 sky130_fd_sc_hd__buf_2 input196 (.A(Tile_X0Y1_E2MID[3]),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(Tile_X0Y1_E2MID[4]),
    .X(net197));
 sky130_fd_sc_hd__buf_2 input198 (.A(Tile_X0Y1_E2MID[5]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input199 (.A(Tile_X0Y1_E2MID[6]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(Tile_X0Y0_E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(Tile_X0Y0_E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input200 (.A(Tile_X0Y1_E2MID[7]),
    .X(net200));
 sky130_fd_sc_hd__buf_4 input201 (.A(Tile_X0Y1_E6END[0]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(Tile_X0Y1_E6END[10]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(Tile_X0Y1_E6END[11]),
    .X(net203));
 sky130_fd_sc_hd__buf_4 input204 (.A(Tile_X0Y1_E6END[1]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(Tile_X0Y1_E6END[2]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(Tile_X0Y1_E6END[3]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(Tile_X0Y1_E6END[4]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(Tile_X0Y1_E6END[5]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(Tile_X0Y1_E6END[6]),
    .X(net209));
 sky130_fd_sc_hd__buf_4 input21 (.A(Tile_X0Y0_E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(Tile_X0Y1_E6END[7]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(Tile_X0Y1_E6END[8]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(Tile_X0Y1_E6END[9]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(Tile_X0Y1_EE4END[0]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(Tile_X0Y1_EE4END[10]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(Tile_X0Y1_EE4END[11]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(Tile_X0Y1_EE4END[12]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(Tile_X0Y1_EE4END[13]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(Tile_X0Y1_EE4END[14]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(Tile_X0Y1_EE4END[15]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(Tile_X0Y0_E6END[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(Tile_X0Y1_EE4END[1]),
    .X(net220));
 sky130_fd_sc_hd__buf_2 input221 (.A(Tile_X0Y1_EE4END[2]),
    .X(net221));
 sky130_fd_sc_hd__buf_1 input222 (.A(Tile_X0Y1_EE4END[3]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(Tile_X0Y1_EE4END[4]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(Tile_X0Y1_EE4END[5]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(Tile_X0Y1_EE4END[6]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(Tile_X0Y1_EE4END[7]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(Tile_X0Y1_EE4END[8]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(Tile_X0Y1_EE4END[9]),
    .X(net228));
 sky130_fd_sc_hd__buf_6 input229 (.A(Tile_X0Y1_FrameData[0]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(Tile_X0Y0_E6END[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_8 input230 (.A(Tile_X0Y1_FrameData[10]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 input231 (.A(Tile_X0Y1_FrameData[11]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_8 input232 (.A(Tile_X0Y1_FrameData[12]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 input233 (.A(Tile_X0Y1_FrameData[13]),
    .X(net233));
 sky130_fd_sc_hd__buf_6 input234 (.A(Tile_X0Y1_FrameData[14]),
    .X(net234));
 sky130_fd_sc_hd__buf_6 input235 (.A(Tile_X0Y1_FrameData[15]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 input236 (.A(Tile_X0Y1_FrameData[16]),
    .X(net236));
 sky130_fd_sc_hd__buf_4 input237 (.A(Tile_X0Y1_FrameData[17]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_8 input238 (.A(Tile_X0Y1_FrameData[18]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_8 input239 (.A(Tile_X0Y1_FrameData[19]),
    .X(net239));
 sky130_fd_sc_hd__buf_4 input24 (.A(Tile_X0Y0_E6END[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 input240 (.A(Tile_X0Y1_FrameData[1]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 input241 (.A(Tile_X0Y1_FrameData[20]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_8 input242 (.A(Tile_X0Y1_FrameData[21]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_8 input243 (.A(Tile_X0Y1_FrameData[22]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_8 input244 (.A(Tile_X0Y1_FrameData[23]),
    .X(net244));
 sky130_fd_sc_hd__buf_4 input245 (.A(Tile_X0Y1_FrameData[24]),
    .X(net245));
 sky130_fd_sc_hd__buf_4 input246 (.A(Tile_X0Y1_FrameData[25]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_8 input247 (.A(Tile_X0Y1_FrameData[26]),
    .X(net247));
 sky130_fd_sc_hd__buf_6 input248 (.A(Tile_X0Y1_FrameData[27]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_8 input249 (.A(Tile_X0Y1_FrameData[28]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(Tile_X0Y0_E6END[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_8 input250 (.A(Tile_X0Y1_FrameData[29]),
    .X(net250));
 sky130_fd_sc_hd__buf_6 input251 (.A(Tile_X0Y1_FrameData[2]),
    .X(net251));
 sky130_fd_sc_hd__buf_6 input252 (.A(Tile_X0Y1_FrameData[30]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 input253 (.A(Tile_X0Y1_FrameData[31]),
    .X(net253));
 sky130_fd_sc_hd__buf_6 input254 (.A(Tile_X0Y1_FrameData[3]),
    .X(net254));
 sky130_fd_sc_hd__buf_6 input255 (.A(Tile_X0Y1_FrameData[4]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 input256 (.A(Tile_X0Y1_FrameData[5]),
    .X(net256));
 sky130_fd_sc_hd__buf_6 input257 (.A(Tile_X0Y1_FrameData[6]),
    .X(net257));
 sky130_fd_sc_hd__buf_6 input258 (.A(Tile_X0Y1_FrameData[7]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 input259 (.A(Tile_X0Y1_FrameData[8]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(Tile_X0Y0_E6END[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_8 input260 (.A(Tile_X0Y1_FrameData[9]),
    .X(net260));
 sky130_fd_sc_hd__buf_8 input261 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net261));
 sky130_fd_sc_hd__buf_8 input262 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net262));
 sky130_fd_sc_hd__buf_8 input263 (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_16 input264 (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 input265 (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 input266 (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 input267 (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 input268 (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 input269 (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(Tile_X0Y0_E6END[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input270 (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 input271 (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(net271));
 sky130_fd_sc_hd__buf_8 input272 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_16 input273 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net273));
 sky130_fd_sc_hd__buf_12 input274 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net274));
 sky130_fd_sc_hd__buf_12 input275 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_16 input276 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net276));
 sky130_fd_sc_hd__buf_8 input277 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net277));
 sky130_fd_sc_hd__buf_8 input278 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net278));
 sky130_fd_sc_hd__buf_8 input279 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(Tile_X0Y0_E6END[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_8 input280 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net280));
 sky130_fd_sc_hd__buf_4 input281 (.A(Tile_X0Y1_N1END[0]),
    .X(net281));
 sky130_fd_sc_hd__buf_4 input282 (.A(Tile_X0Y1_N1END[1]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 input283 (.A(Tile_X0Y1_N1END[2]),
    .X(net283));
 sky130_fd_sc_hd__buf_4 input284 (.A(Tile_X0Y1_N1END[3]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 input285 (.A(Tile_X0Y1_N2END[0]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 input286 (.A(Tile_X0Y1_N2END[1]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 input287 (.A(Tile_X0Y1_N2END[2]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 input288 (.A(Tile_X0Y1_N2END[3]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 input289 (.A(Tile_X0Y1_N2END[4]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(Tile_X0Y0_E6END[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input290 (.A(Tile_X0Y1_N2END[5]),
    .X(net290));
 sky130_fd_sc_hd__buf_2 input291 (.A(Tile_X0Y1_N2END[6]),
    .X(net291));
 sky130_fd_sc_hd__buf_2 input292 (.A(Tile_X0Y1_N2END[7]),
    .X(net292));
 sky130_fd_sc_hd__buf_2 input293 (.A(Tile_X0Y1_N2MID[0]),
    .X(net293));
 sky130_fd_sc_hd__buf_2 input294 (.A(Tile_X0Y1_N2MID[1]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 input295 (.A(Tile_X0Y1_N2MID[2]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 input296 (.A(Tile_X0Y1_N2MID[3]),
    .X(net296));
 sky130_fd_sc_hd__buf_2 input297 (.A(Tile_X0Y1_N2MID[4]),
    .X(net297));
 sky130_fd_sc_hd__buf_2 input298 (.A(Tile_X0Y1_N2MID[5]),
    .X(net298));
 sky130_fd_sc_hd__buf_4 input299 (.A(Tile_X0Y1_N2MID[6]),
    .X(net299));
 sky130_fd_sc_hd__buf_4 input3 (.A(Tile_X0Y0_E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(Tile_X0Y0_E6END[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input300 (.A(Tile_X0Y1_N2MID[7]),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 input301 (.A(Tile_X0Y1_N4END[0]),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 input302 (.A(Tile_X0Y1_N4END[10]),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 input303 (.A(Tile_X0Y1_N4END[11]),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 input304 (.A(Tile_X0Y1_N4END[12]),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 input305 (.A(Tile_X0Y1_N4END[13]),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 input306 (.A(Tile_X0Y1_N4END[14]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 input307 (.A(Tile_X0Y1_N4END[15]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 input308 (.A(Tile_X0Y1_N4END[1]),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 input309 (.A(Tile_X0Y1_N4END[2]),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(Tile_X0Y0_E6END[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input310 (.A(Tile_X0Y1_N4END[3]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(Tile_X0Y1_N4END[4]),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 input312 (.A(Tile_X0Y1_N4END[5]),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 input313 (.A(Tile_X0Y1_N4END[6]),
    .X(net313));
 sky130_fd_sc_hd__buf_2 input314 (.A(Tile_X0Y1_N4END[7]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 input315 (.A(Tile_X0Y1_N4END[8]),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 input316 (.A(Tile_X0Y1_N4END[9]),
    .X(net316));
 sky130_fd_sc_hd__buf_1 input317 (.A(Tile_X0Y1_NN4END[0]),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 input318 (.A(Tile_X0Y1_NN4END[10]),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 input319 (.A(Tile_X0Y1_NN4END[11]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(Tile_X0Y0_E6END[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input320 (.A(Tile_X0Y1_NN4END[12]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 input321 (.A(Tile_X0Y1_NN4END[13]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 input322 (.A(Tile_X0Y1_NN4END[14]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 input323 (.A(Tile_X0Y1_NN4END[15]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 input324 (.A(Tile_X0Y1_NN4END[1]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 input325 (.A(Tile_X0Y1_NN4END[2]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 input326 (.A(Tile_X0Y1_NN4END[3]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 input327 (.A(Tile_X0Y1_NN4END[4]),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 input328 (.A(Tile_X0Y1_NN4END[5]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 input329 (.A(Tile_X0Y1_NN4END[6]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(Tile_X0Y0_EE4END[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input330 (.A(Tile_X0Y1_NN4END[7]),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 input331 (.A(Tile_X0Y1_NN4END[8]),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 input332 (.A(Tile_X0Y1_NN4END[9]),
    .X(net332));
 sky130_fd_sc_hd__buf_12 input333 (.A(Tile_X0Y1_UserCLK),
    .X(net333));
 sky130_fd_sc_hd__buf_4 input334 (.A(Tile_X0Y1_W1END[0]),
    .X(net334));
 sky130_fd_sc_hd__buf_4 input335 (.A(Tile_X0Y1_W1END[1]),
    .X(net335));
 sky130_fd_sc_hd__buf_4 input336 (.A(Tile_X0Y1_W1END[2]),
    .X(net336));
 sky130_fd_sc_hd__buf_4 input337 (.A(Tile_X0Y1_W1END[3]),
    .X(net337));
 sky130_fd_sc_hd__buf_2 input338 (.A(Tile_X0Y1_W2END[0]),
    .X(net338));
 sky130_fd_sc_hd__buf_2 input339 (.A(Tile_X0Y1_W2END[1]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(Tile_X0Y0_EE4END[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input340 (.A(Tile_X0Y1_W2END[2]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 input341 (.A(Tile_X0Y1_W2END[3]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 input342 (.A(Tile_X0Y1_W2END[4]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 input343 (.A(Tile_X0Y1_W2END[5]),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 input344 (.A(Tile_X0Y1_W2END[6]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 input345 (.A(Tile_X0Y1_W2END[7]),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 input346 (.A(Tile_X0Y1_W2MID[0]),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 input347 (.A(Tile_X0Y1_W2MID[1]),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_4 input348 (.A(Tile_X0Y1_W2MID[2]),
    .X(net348));
 sky130_fd_sc_hd__buf_2 input349 (.A(Tile_X0Y1_W2MID[3]),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(Tile_X0Y0_EE4END[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input350 (.A(Tile_X0Y1_W2MID[4]),
    .X(net350));
 sky130_fd_sc_hd__buf_2 input351 (.A(Tile_X0Y1_W2MID[5]),
    .X(net351));
 sky130_fd_sc_hd__buf_4 input352 (.A(Tile_X0Y1_W2MID[6]),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_4 input353 (.A(Tile_X0Y1_W2MID[7]),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 input354 (.A(Tile_X0Y1_W6END[0]),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 input355 (.A(Tile_X0Y1_W6END[10]),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 input356 (.A(Tile_X0Y1_W6END[11]),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 input357 (.A(Tile_X0Y1_W6END[1]),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 input358 (.A(Tile_X0Y1_W6END[2]),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 input359 (.A(Tile_X0Y1_W6END[3]),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(Tile_X0Y0_EE4END[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input360 (.A(Tile_X0Y1_W6END[4]),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 input361 (.A(Tile_X0Y1_W6END[5]),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 input362 (.A(Tile_X0Y1_W6END[6]),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 input363 (.A(Tile_X0Y1_W6END[7]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 input364 (.A(Tile_X0Y1_W6END[8]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 input365 (.A(Tile_X0Y1_W6END[9]),
    .X(net365));
 sky130_fd_sc_hd__buf_2 input366 (.A(Tile_X0Y1_WW4END[0]),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 input367 (.A(Tile_X0Y1_WW4END[10]),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 input368 (.A(Tile_X0Y1_WW4END[11]),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 input369 (.A(Tile_X0Y1_WW4END[12]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(Tile_X0Y0_EE4END[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input370 (.A(Tile_X0Y1_WW4END[13]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 input371 (.A(Tile_X0Y1_WW4END[14]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 input372 (.A(Tile_X0Y1_WW4END[15]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 input373 (.A(Tile_X0Y1_WW4END[1]),
    .X(net373));
 sky130_fd_sc_hd__buf_2 input374 (.A(Tile_X0Y1_WW4END[2]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 input375 (.A(Tile_X0Y1_WW4END[3]),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 input376 (.A(Tile_X0Y1_WW4END[4]),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 input377 (.A(Tile_X0Y1_WW4END[5]),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 input378 (.A(Tile_X0Y1_WW4END[6]),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 input379 (.A(Tile_X0Y1_WW4END[7]),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(Tile_X0Y0_EE4END[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input380 (.A(Tile_X0Y1_WW4END[8]),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 input381 (.A(Tile_X0Y1_WW4END[9]),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(Tile_X0Y0_EE4END[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(Tile_X0Y0_E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(Tile_X0Y0_EE4END[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(Tile_X0Y0_EE4END[2]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(Tile_X0Y0_EE4END[3]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(Tile_X0Y0_EE4END[4]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(Tile_X0Y0_EE4END[5]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(Tile_X0Y0_EE4END[6]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(Tile_X0Y0_EE4END[7]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(Tile_X0Y0_EE4END[8]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(Tile_X0Y0_EE4END[9]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(Tile_X0Y0_FrameData[0]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(Tile_X0Y0_E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(Tile_X0Y0_FrameData[10]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(Tile_X0Y0_FrameData[11]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_8 input52 (.A(Tile_X0Y0_FrameData[12]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 input53 (.A(Tile_X0Y0_FrameData[13]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 input54 (.A(Tile_X0Y0_FrameData[14]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 input55 (.A(Tile_X0Y0_FrameData[15]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 input56 (.A(Tile_X0Y0_FrameData[16]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 input57 (.A(Tile_X0Y0_FrameData[17]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 input58 (.A(Tile_X0Y0_FrameData[18]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(Tile_X0Y0_FrameData[19]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(Tile_X0Y0_E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input60 (.A(Tile_X0Y0_FrameData[1]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 input61 (.A(Tile_X0Y0_FrameData[20]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 input62 (.A(Tile_X0Y0_FrameData[21]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(Tile_X0Y0_FrameData[22]),
    .X(net63));
 sky130_fd_sc_hd__buf_6 input64 (.A(Tile_X0Y0_FrameData[23]),
    .X(net64));
 sky130_fd_sc_hd__buf_6 input65 (.A(Tile_X0Y0_FrameData[24]),
    .X(net65));
 sky130_fd_sc_hd__buf_6 input66 (.A(Tile_X0Y0_FrameData[25]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(Tile_X0Y0_FrameData[26]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 input68 (.A(Tile_X0Y0_FrameData[27]),
    .X(net68));
 sky130_fd_sc_hd__buf_6 input69 (.A(Tile_X0Y0_FrameData[28]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(Tile_X0Y0_E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input70 (.A(Tile_X0Y0_FrameData[29]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 input71 (.A(Tile_X0Y0_FrameData[2]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 input72 (.A(Tile_X0Y0_FrameData[30]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 input73 (.A(Tile_X0Y0_FrameData[31]),
    .X(net73));
 sky130_fd_sc_hd__buf_6 input74 (.A(Tile_X0Y0_FrameData[3]),
    .X(net74));
 sky130_fd_sc_hd__buf_6 input75 (.A(Tile_X0Y0_FrameData[4]),
    .X(net75));
 sky130_fd_sc_hd__buf_6 input76 (.A(Tile_X0Y0_FrameData[5]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 input77 (.A(Tile_X0Y0_FrameData[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 input78 (.A(Tile_X0Y0_FrameData[7]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(Tile_X0Y0_FrameData[8]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(Tile_X0Y0_E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(Tile_X0Y0_FrameData[9]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(Tile_X0Y0_S1END[0]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(Tile_X0Y0_S1END[1]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(Tile_X0Y0_S1END[2]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(Tile_X0Y0_S1END[3]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(Tile_X0Y0_S2END[0]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(Tile_X0Y0_S2END[1]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(Tile_X0Y0_S2END[2]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(Tile_X0Y0_S2END[3]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(Tile_X0Y0_S2END[4]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(Tile_X0Y0_E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input90 (.A(Tile_X0Y0_S2END[5]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(Tile_X0Y0_S2END[6]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(Tile_X0Y0_S2END[7]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(Tile_X0Y0_S2MID[0]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(Tile_X0Y0_S2MID[1]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 input95 (.A(Tile_X0Y0_S2MID[2]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 input96 (.A(Tile_X0Y0_S2MID[3]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 input97 (.A(Tile_X0Y0_S2MID[4]),
    .X(net97));
 sky130_fd_sc_hd__buf_4 input98 (.A(Tile_X0Y0_S2MID[5]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(Tile_X0Y0_S2MID[6]),
    .X(net99));
 sky130_fd_sc_hd__buf_12 max_cap763 (.A(\Tile_X0Y1_DSP_bot/Q6 ),
    .X(net763));
 sky130_fd_sc_hd__buf_6 max_cap764 (.A(\Tile_X0Y1_DSP_bot/Q1 ),
    .X(net764));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(Tile_X0Y0_E1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .X(Tile_X0Y0_E1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(Tile_X0Y0_E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .X(Tile_X0Y0_E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(Tile_X0Y0_E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .X(Tile_X0Y0_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(Tile_X0Y0_E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .X(Tile_X0Y0_E2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .X(Tile_X0Y0_E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output391 (.A(net391),
    .X(Tile_X0Y0_E2BEG[5]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(Tile_X0Y0_E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output393 (.A(net393),
    .X(Tile_X0Y0_E2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output394 (.A(net394),
    .X(Tile_X0Y0_E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output395 (.A(net395),
    .X(Tile_X0Y0_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .X(Tile_X0Y0_E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output397 (.A(net397),
    .X(Tile_X0Y0_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net398),
    .X(Tile_X0Y0_E2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output399 (.A(net399),
    .X(Tile_X0Y0_E2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output400 (.A(net400),
    .X(Tile_X0Y0_E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output401 (.A(net401),
    .X(Tile_X0Y0_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net402),
    .X(Tile_X0Y0_E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net403),
    .X(Tile_X0Y0_E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output404 (.A(net404),
    .X(Tile_X0Y0_E6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output405 (.A(net405),
    .X(Tile_X0Y0_E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output406 (.A(net406),
    .X(Tile_X0Y0_E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output407 (.A(net407),
    .X(Tile_X0Y0_E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .X(Tile_X0Y0_E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output409 (.A(net409),
    .X(Tile_X0Y0_E6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output410 (.A(net410),
    .X(Tile_X0Y0_E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output411 (.A(net411),
    .X(Tile_X0Y0_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(Tile_X0Y0_E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output413 (.A(net413),
    .X(Tile_X0Y0_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .X(Tile_X0Y0_EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(Tile_X0Y0_EE4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output416 (.A(net416),
    .X(Tile_X0Y0_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .X(Tile_X0Y0_EE4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output418 (.A(net418),
    .X(Tile_X0Y0_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .X(Tile_X0Y0_EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output420 (.A(net420),
    .X(Tile_X0Y0_EE4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output421 (.A(net421),
    .X(Tile_X0Y0_EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output422 (.A(net422),
    .X(Tile_X0Y0_EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output423 (.A(net423),
    .X(Tile_X0Y0_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net424),
    .X(Tile_X0Y0_EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output425 (.A(net425),
    .X(Tile_X0Y0_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .X(Tile_X0Y0_EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output427 (.A(net427),
    .X(Tile_X0Y0_EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output428 (.A(net428),
    .X(Tile_X0Y0_EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output429 (.A(net429),
    .X(Tile_X0Y0_EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output430 (.A(net430),
    .X(Tile_X0Y0_FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output431 (.A(net431),
    .X(Tile_X0Y0_FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output432 (.A(net432),
    .X(Tile_X0Y0_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .X(Tile_X0Y0_FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output434 (.A(net434),
    .X(Tile_X0Y0_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net435),
    .X(Tile_X0Y0_FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output436 (.A(net436),
    .X(Tile_X0Y0_FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output437 (.A(net437),
    .X(Tile_X0Y0_FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output438 (.A(net438),
    .X(Tile_X0Y0_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .X(Tile_X0Y0_FrameData_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output440 (.A(net440),
    .X(Tile_X0Y0_FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output441 (.A(net441),
    .X(Tile_X0Y0_FrameData_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output442 (.A(net442),
    .X(Tile_X0Y0_FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output443 (.A(net443),
    .X(Tile_X0Y0_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net444),
    .X(Tile_X0Y0_FrameData_O[22]));
 sky130_fd_sc_hd__clkbuf_4 output445 (.A(net445),
    .X(Tile_X0Y0_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output446 (.A(net446),
    .X(Tile_X0Y0_FrameData_O[24]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .X(Tile_X0Y0_FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output448 (.A(net448),
    .X(Tile_X0Y0_FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output449 (.A(net449),
    .X(Tile_X0Y0_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .X(Tile_X0Y0_FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output451 (.A(net451),
    .X(Tile_X0Y0_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .X(Tile_X0Y0_FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output453 (.A(net453),
    .X(Tile_X0Y0_FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output454 (.A(net454),
    .X(Tile_X0Y0_FrameData_O[31]));
 sky130_fd_sc_hd__clkbuf_4 output455 (.A(net455),
    .X(Tile_X0Y0_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .X(Tile_X0Y0_FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output457 (.A(net457),
    .X(Tile_X0Y0_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net458),
    .X(Tile_X0Y0_FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output459 (.A(net459),
    .X(Tile_X0Y0_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .X(Tile_X0Y0_FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output461 (.A(net461),
    .X(Tile_X0Y0_FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output462 (.A(net462),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output463 (.A(net463),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output464 (.A(net464),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output467 (.A(net467),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output468 (.A(net468),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output469 (.A(net469),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output470 (.A(net470),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output471 (.A(net471),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output472 (.A(net472),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output473 (.A(net473),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net474),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output475 (.A(net475),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output476 (.A(net476),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output477 (.A(net477),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output478 (.A(net478),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output479 (.A(net479),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output480 (.A(net480),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output481 (.A(net481),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output482 (.A(net482),
    .X(Tile_X0Y0_N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output483 (.A(net483),
    .X(Tile_X0Y0_N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output484 (.A(net484),
    .X(Tile_X0Y0_N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output485 (.A(net485),
    .X(Tile_X0Y0_N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .X(Tile_X0Y0_N2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output487 (.A(net487),
    .X(Tile_X0Y0_N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output488 (.A(net488),
    .X(Tile_X0Y0_N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output489 (.A(net489),
    .X(Tile_X0Y0_N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net490),
    .X(Tile_X0Y0_N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output491 (.A(net491),
    .X(Tile_X0Y0_N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net492),
    .X(Tile_X0Y0_N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output493 (.A(net493),
    .X(Tile_X0Y0_N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output494 (.A(net494),
    .X(Tile_X0Y0_N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net495),
    .X(Tile_X0Y0_N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net496),
    .X(Tile_X0Y0_N2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output497 (.A(net497),
    .X(Tile_X0Y0_N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net498),
    .X(Tile_X0Y0_N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output499 (.A(net499),
    .X(Tile_X0Y0_N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .X(Tile_X0Y0_N2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output501 (.A(net501),
    .X(Tile_X0Y0_N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net502),
    .X(Tile_X0Y0_N4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output503 (.A(net503),
    .X(Tile_X0Y0_N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output504 (.A(net504),
    .X(Tile_X0Y0_N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output505 (.A(net505),
    .X(Tile_X0Y0_N4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output506 (.A(net506),
    .X(Tile_X0Y0_N4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output507 (.A(net507),
    .X(Tile_X0Y0_N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output508 (.A(net508),
    .X(Tile_X0Y0_N4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output509 (.A(net509),
    .X(Tile_X0Y0_N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output510 (.A(net510),
    .X(Tile_X0Y0_N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output511 (.A(net511),
    .X(Tile_X0Y0_N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output512 (.A(net512),
    .X(Tile_X0Y0_N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output513 (.A(net513),
    .X(Tile_X0Y0_N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output514 (.A(net514),
    .X(Tile_X0Y0_N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output515 (.A(net515),
    .X(Tile_X0Y0_N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output516 (.A(net516),
    .X(Tile_X0Y0_N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output517 (.A(net517),
    .X(Tile_X0Y0_N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output518 (.A(net518),
    .X(Tile_X0Y0_NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output519 (.A(net519),
    .X(Tile_X0Y0_NN4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output520 (.A(net520),
    .X(Tile_X0Y0_NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output521 (.A(net521),
    .X(Tile_X0Y0_NN4BEG[12]));
 sky130_fd_sc_hd__buf_2 output522 (.A(net522),
    .X(Tile_X0Y0_NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output523 (.A(net523),
    .X(Tile_X0Y0_NN4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output524 (.A(net524),
    .X(Tile_X0Y0_NN4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output525 (.A(net525),
    .X(Tile_X0Y0_NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output526 (.A(net526),
    .X(Tile_X0Y0_NN4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output527 (.A(net527),
    .X(Tile_X0Y0_NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output528 (.A(net528),
    .X(Tile_X0Y0_NN4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output529 (.A(net529),
    .X(Tile_X0Y0_NN4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output530 (.A(net530),
    .X(Tile_X0Y0_NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output531 (.A(net531),
    .X(Tile_X0Y0_NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output532 (.A(net532),
    .X(Tile_X0Y0_NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output533 (.A(net533),
    .X(Tile_X0Y0_NN4BEG[9]));
 sky130_fd_sc_hd__buf_2 output534 (.A(net534),
    .X(Tile_X0Y0_UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output535 (.A(net535),
    .X(Tile_X0Y0_W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output536 (.A(net536),
    .X(Tile_X0Y0_W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output537 (.A(net537),
    .X(Tile_X0Y0_W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output538 (.A(net538),
    .X(Tile_X0Y0_W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output539 (.A(net539),
    .X(Tile_X0Y0_W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output540 (.A(net540),
    .X(Tile_X0Y0_W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output541 (.A(net541),
    .X(Tile_X0Y0_W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output542 (.A(net542),
    .X(Tile_X0Y0_W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output543 (.A(net543),
    .X(Tile_X0Y0_W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output544 (.A(net544),
    .X(Tile_X0Y0_W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output545 (.A(net545),
    .X(Tile_X0Y0_W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output546 (.A(net546),
    .X(Tile_X0Y0_W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output547 (.A(net547),
    .X(Tile_X0Y0_W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output548 (.A(net548),
    .X(Tile_X0Y0_W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output549 (.A(net549),
    .X(Tile_X0Y0_W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output550 (.A(net550),
    .X(Tile_X0Y0_W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output551 (.A(net551),
    .X(Tile_X0Y0_W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output552 (.A(net552),
    .X(Tile_X0Y0_W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output553 (.A(net553),
    .X(Tile_X0Y0_W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output554 (.A(net554),
    .X(Tile_X0Y0_W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output555 (.A(net555),
    .X(Tile_X0Y0_W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output556 (.A(net556),
    .X(Tile_X0Y0_W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output557 (.A(net557),
    .X(Tile_X0Y0_W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output558 (.A(net558),
    .X(Tile_X0Y0_W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output559 (.A(net559),
    .X(Tile_X0Y0_W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output560 (.A(net560),
    .X(Tile_X0Y0_W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output561 (.A(net561),
    .X(Tile_X0Y0_W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output562 (.A(net562),
    .X(Tile_X0Y0_W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output563 (.A(net563),
    .X(Tile_X0Y0_W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output564 (.A(net564),
    .X(Tile_X0Y0_W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output565 (.A(net565),
    .X(Tile_X0Y0_W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output566 (.A(net566),
    .X(Tile_X0Y0_W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output567 (.A(net567),
    .X(Tile_X0Y0_WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output568 (.A(net568),
    .X(Tile_X0Y0_WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output569 (.A(net569),
    .X(Tile_X0Y0_WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output570 (.A(net570),
    .X(Tile_X0Y0_WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output571 (.A(net571),
    .X(Tile_X0Y0_WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output572 (.A(net572),
    .X(Tile_X0Y0_WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output573 (.A(net573),
    .X(Tile_X0Y0_WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output574 (.A(net574),
    .X(Tile_X0Y0_WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output575 (.A(net575),
    .X(Tile_X0Y0_WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output576 (.A(net576),
    .X(Tile_X0Y0_WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output577 (.A(net577),
    .X(Tile_X0Y0_WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output578 (.A(net578),
    .X(Tile_X0Y0_WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output579 (.A(net579),
    .X(Tile_X0Y0_WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output580 (.A(net580),
    .X(Tile_X0Y0_WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output581 (.A(net581),
    .X(Tile_X0Y0_WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output582 (.A(net582),
    .X(Tile_X0Y0_WW4BEG[9]));
 sky130_fd_sc_hd__buf_2 output583 (.A(net583),
    .X(Tile_X0Y1_E1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output584 (.A(net584),
    .X(Tile_X0Y1_E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output585 (.A(net585),
    .X(Tile_X0Y1_E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output586 (.A(net586),
    .X(Tile_X0Y1_E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output587 (.A(net587),
    .X(Tile_X0Y1_E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output588 (.A(net588),
    .X(Tile_X0Y1_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output589 (.A(net589),
    .X(Tile_X0Y1_E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output590 (.A(net590),
    .X(Tile_X0Y1_E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output591 (.A(net591),
    .X(Tile_X0Y1_E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output592 (.A(net592),
    .X(Tile_X0Y1_E2BEG[5]));
 sky130_fd_sc_hd__buf_2 output593 (.A(net593),
    .X(Tile_X0Y1_E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output594 (.A(net594),
    .X(Tile_X0Y1_E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output595 (.A(net595),
    .X(Tile_X0Y1_E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output596 (.A(net596),
    .X(Tile_X0Y1_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output597 (.A(net597),
    .X(Tile_X0Y1_E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output598 (.A(net598),
    .X(Tile_X0Y1_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output599 (.A(net599),
    .X(Tile_X0Y1_E2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output600 (.A(net600),
    .X(Tile_X0Y1_E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output601 (.A(net601),
    .X(Tile_X0Y1_E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output602 (.A(net602),
    .X(Tile_X0Y1_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output603 (.A(net603),
    .X(Tile_X0Y1_E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output604 (.A(net604),
    .X(Tile_X0Y1_E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output605 (.A(net605),
    .X(Tile_X0Y1_E6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output606 (.A(net606),
    .X(Tile_X0Y1_E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output607 (.A(net607),
    .X(Tile_X0Y1_E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output608 (.A(net608),
    .X(Tile_X0Y1_E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output609 (.A(net609),
    .X(Tile_X0Y1_E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output610 (.A(net610),
    .X(Tile_X0Y1_E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output611 (.A(net611),
    .X(Tile_X0Y1_E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output612 (.A(net612),
    .X(Tile_X0Y1_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output613 (.A(net613),
    .X(Tile_X0Y1_E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output614 (.A(net614),
    .X(Tile_X0Y1_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output615 (.A(net615),
    .X(Tile_X0Y1_EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output616 (.A(net616),
    .X(Tile_X0Y1_EE4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output617 (.A(net617),
    .X(Tile_X0Y1_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output618 (.A(net618),
    .X(Tile_X0Y1_EE4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output619 (.A(net619),
    .X(Tile_X0Y1_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output620 (.A(net620),
    .X(Tile_X0Y1_EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output621 (.A(net621),
    .X(Tile_X0Y1_EE4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output622 (.A(net622),
    .X(Tile_X0Y1_EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output623 (.A(net623),
    .X(Tile_X0Y1_EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output624 (.A(net624),
    .X(Tile_X0Y1_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output625 (.A(net625),
    .X(Tile_X0Y1_EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output626 (.A(net626),
    .X(Tile_X0Y1_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output627 (.A(net627),
    .X(Tile_X0Y1_EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output628 (.A(net628),
    .X(Tile_X0Y1_EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output629 (.A(net629),
    .X(Tile_X0Y1_EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output630 (.A(net630),
    .X(Tile_X0Y1_EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output631 (.A(net631),
    .X(Tile_X0Y1_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output632 (.A(net632),
    .X(Tile_X0Y1_FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output633 (.A(net633),
    .X(Tile_X0Y1_FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output634 (.A(net634),
    .X(Tile_X0Y1_FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output635 (.A(net635),
    .X(Tile_X0Y1_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output636 (.A(net636),
    .X(Tile_X0Y1_FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output637 (.A(net637),
    .X(Tile_X0Y1_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output638 (.A(net638),
    .X(Tile_X0Y1_FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output639 (.A(net639),
    .X(Tile_X0Y1_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output640 (.A(net640),
    .X(Tile_X0Y1_FrameData_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output641 (.A(net641),
    .X(Tile_X0Y1_FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output642 (.A(net642),
    .X(Tile_X0Y1_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output643 (.A(net643),
    .X(Tile_X0Y1_FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output644 (.A(net644),
    .X(Tile_X0Y1_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output645 (.A(net645),
    .X(Tile_X0Y1_FrameData_O[22]));
 sky130_fd_sc_hd__clkbuf_4 output646 (.A(net646),
    .X(Tile_X0Y1_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output647 (.A(net647),
    .X(Tile_X0Y1_FrameData_O[24]));
 sky130_fd_sc_hd__clkbuf_4 output648 (.A(net648),
    .X(Tile_X0Y1_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output649 (.A(net649),
    .X(Tile_X0Y1_FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output650 (.A(net650),
    .X(Tile_X0Y1_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output651 (.A(net651),
    .X(Tile_X0Y1_FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output652 (.A(net652),
    .X(Tile_X0Y1_FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output653 (.A(net653),
    .X(Tile_X0Y1_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output654 (.A(net654),
    .X(Tile_X0Y1_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output655 (.A(net655),
    .X(Tile_X0Y1_FrameData_O[31]));
 sky130_fd_sc_hd__clkbuf_4 output656 (.A(net656),
    .X(Tile_X0Y1_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output657 (.A(net657),
    .X(Tile_X0Y1_FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output658 (.A(net658),
    .X(Tile_X0Y1_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output659 (.A(net659),
    .X(Tile_X0Y1_FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output660 (.A(net660),
    .X(Tile_X0Y1_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output661 (.A(net661),
    .X(Tile_X0Y1_FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output662 (.A(net662),
    .X(Tile_X0Y1_FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output663 (.A(net663),
    .X(Tile_X0Y1_S1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output664 (.A(net664),
    .X(Tile_X0Y1_S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output665 (.A(net665),
    .X(Tile_X0Y1_S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output666 (.A(net666),
    .X(Tile_X0Y1_S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output667 (.A(net667),
    .X(Tile_X0Y1_S2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output668 (.A(net668),
    .X(Tile_X0Y1_S2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output669 (.A(net669),
    .X(Tile_X0Y1_S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output670 (.A(net670),
    .X(Tile_X0Y1_S2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output671 (.A(net671),
    .X(Tile_X0Y1_S2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output672 (.A(net672),
    .X(Tile_X0Y1_S2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output673 (.A(net673),
    .X(Tile_X0Y1_S2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output674 (.A(net674),
    .X(Tile_X0Y1_S2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output675 (.A(net675),
    .X(Tile_X0Y1_S2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output676 (.A(net676),
    .X(Tile_X0Y1_S2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output677 (.A(net677),
    .X(Tile_X0Y1_S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output678 (.A(net678),
    .X(Tile_X0Y1_S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output679 (.A(net679),
    .X(Tile_X0Y1_S2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output680 (.A(net680),
    .X(Tile_X0Y1_S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output681 (.A(net681),
    .X(Tile_X0Y1_S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output682 (.A(net682),
    .X(Tile_X0Y1_S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output683 (.A(net683),
    .X(Tile_X0Y1_S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output684 (.A(net684),
    .X(Tile_X0Y1_S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output685 (.A(net685),
    .X(Tile_X0Y1_S4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output686 (.A(net686),
    .X(Tile_X0Y1_S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output687 (.A(net687),
    .X(Tile_X0Y1_S4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output688 (.A(net688),
    .X(Tile_X0Y1_S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output689 (.A(net689),
    .X(Tile_X0Y1_S4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output690 (.A(net690),
    .X(Tile_X0Y1_S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output691 (.A(net691),
    .X(Tile_X0Y1_S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output692 (.A(net692),
    .X(Tile_X0Y1_S4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output693 (.A(net693),
    .X(Tile_X0Y1_S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output694 (.A(net694),
    .X(Tile_X0Y1_S4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output695 (.A(net695),
    .X(Tile_X0Y1_S4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output696 (.A(net696),
    .X(Tile_X0Y1_S4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output697 (.A(net697),
    .X(Tile_X0Y1_S4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output698 (.A(net698),
    .X(Tile_X0Y1_S4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output699 (.A(net699),
    .X(Tile_X0Y1_SS4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output700 (.A(net700),
    .X(Tile_X0Y1_SS4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output701 (.A(net701),
    .X(Tile_X0Y1_SS4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output702 (.A(net702),
    .X(Tile_X0Y1_SS4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output703 (.A(net703),
    .X(Tile_X0Y1_SS4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output704 (.A(net704),
    .X(Tile_X0Y1_SS4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output705 (.A(net705),
    .X(Tile_X0Y1_SS4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output706 (.A(net706),
    .X(Tile_X0Y1_SS4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output707 (.A(net707),
    .X(Tile_X0Y1_SS4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output708 (.A(net708),
    .X(Tile_X0Y1_SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output709 (.A(net709),
    .X(Tile_X0Y1_SS4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output710 (.A(net710),
    .X(Tile_X0Y1_SS4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output711 (.A(net711),
    .X(Tile_X0Y1_SS4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output712 (.A(net712),
    .X(Tile_X0Y1_SS4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output713 (.A(net713),
    .X(Tile_X0Y1_SS4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output714 (.A(net714),
    .X(Tile_X0Y1_SS4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output715 (.A(net715),
    .X(Tile_X0Y1_W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output716 (.A(net716),
    .X(Tile_X0Y1_W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output717 (.A(net717),
    .X(Tile_X0Y1_W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output718 (.A(net718),
    .X(Tile_X0Y1_W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output719 (.A(net719),
    .X(Tile_X0Y1_W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output720 (.A(net720),
    .X(Tile_X0Y1_W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output721 (.A(net721),
    .X(Tile_X0Y1_W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output722 (.A(net722),
    .X(Tile_X0Y1_W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output723 (.A(net723),
    .X(Tile_X0Y1_W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output724 (.A(net724),
    .X(Tile_X0Y1_W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output725 (.A(net725),
    .X(Tile_X0Y1_W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output726 (.A(net726),
    .X(Tile_X0Y1_W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output727 (.A(net727),
    .X(Tile_X0Y1_W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output728 (.A(net728),
    .X(Tile_X0Y1_W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output729 (.A(net729),
    .X(Tile_X0Y1_W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output730 (.A(net730),
    .X(Tile_X0Y1_W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output731 (.A(net731),
    .X(Tile_X0Y1_W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output732 (.A(net732),
    .X(Tile_X0Y1_W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output733 (.A(net733),
    .X(Tile_X0Y1_W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output734 (.A(net734),
    .X(Tile_X0Y1_W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output735 (.A(net735),
    .X(Tile_X0Y1_W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output736 (.A(net736),
    .X(Tile_X0Y1_W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output737 (.A(net737),
    .X(Tile_X0Y1_W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output738 (.A(net738),
    .X(Tile_X0Y1_W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output739 (.A(net739),
    .X(Tile_X0Y1_W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output740 (.A(net740),
    .X(Tile_X0Y1_W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output741 (.A(net741),
    .X(Tile_X0Y1_W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output742 (.A(net742),
    .X(Tile_X0Y1_W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output743 (.A(net743),
    .X(Tile_X0Y1_W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output744 (.A(net744),
    .X(Tile_X0Y1_W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output745 (.A(net745),
    .X(Tile_X0Y1_W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output746 (.A(net746),
    .X(Tile_X0Y1_W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output747 (.A(net747),
    .X(Tile_X0Y1_WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output748 (.A(net748),
    .X(Tile_X0Y1_WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output749 (.A(net749),
    .X(Tile_X0Y1_WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output750 (.A(net750),
    .X(Tile_X0Y1_WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output751 (.A(net751),
    .X(Tile_X0Y1_WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output752 (.A(net752),
    .X(Tile_X0Y1_WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output753 (.A(net753),
    .X(Tile_X0Y1_WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output754 (.A(net754),
    .X(Tile_X0Y1_WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output755 (.A(net755),
    .X(Tile_X0Y1_WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output756 (.A(net756),
    .X(Tile_X0Y1_WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output757 (.A(net757),
    .X(Tile_X0Y1_WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output758 (.A(net758),
    .X(Tile_X0Y1_WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output759 (.A(net759),
    .X(Tile_X0Y1_WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output760 (.A(net760),
    .X(Tile_X0Y1_WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output761 (.A(net761),
    .X(Tile_X0Y1_WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output762 (.A(net762),
    .X(Tile_X0Y1_WW4BEG[9]));
endmodule

